* E:\smaslan\LV_prog\open-z-bridge-master\sim\LiB_brg_2x4T_twax.asc
XZ1 N046 N050 N047 N051 STDCOAX Rp={Rp1} Lp={Lp1} Rpg={Rp1r} Lpg={Lp1r} kp={kpo1} Cps={Cp1s} Rps={Rp1s} Rc={Rc1} Lc={Lc1} Rcg={Rc1r} Lcg={Lc1r} kc={kco1} Ccs={Cc1s} Rcs={Rc1s} Rs={R1} Ls={L1}
* <component=coax_joint>Rs=Rc3h Ls=Lc3h RsG=Rc3g LsG=Lc3g Cp=Cc3sh Rp=Rc3sh k=kc3 Rch=Rc3ch </component>
.param Rs2_COAXCAB01={0.5*Rc3h} Ls2_COAXCAB01={0.5*Lc3h} RsG2_COAXCAB01={0.5*Rc3g} LsG2_COAXCAB01={0.5*Lc3g} 
R1COAXCAB01 N038 n001COAXCAB01 {Rs2_COAXCAB01} 
L1COAXCAB01 n001COAXCAB01 n002COAXCAB01 {Ls2_COAXCAB01} 
L2COAXCAB01 n002COAXCAB01 n003COAXCAB01 {Ls2_COAXCAB01} 
R2COAXCAB01 n003COAXCAB01 n007COAXCAB01 {Rs2_COAXCAB01} 
K1COAXCAB01 L1COAXCAB01 L3COAXCAB01 {kc3} 
R3COAXCAB01 N029 n004COAXCAB01 {RsG2_COAXCAB01} 
L3COAXCAB01 n004COAXCAB01 n005COAXCAB01 {LsG2_COAXCAB01} 
L4COAXCAB01 n005COAXCAB01 n006COAXCAB01 {LsG2_COAXCAB01} 
R4COAXCAB01 n006COAXCAB01 n009COAXCAB01 {RsG2_COAXCAB01} 
K2COAXCAB01 L2COAXCAB01 L4COAXCAB01 {kc3} 
C1COAXCAB01 n002COAXCAB01 n005COAXCAB01 {Cc3sh} 
R5COAXCAB01 n002COAXCAB01 n005COAXCAB01 {Rc3sh} 
R6COAXCAB01 n007COAXCAB01 n008COAXCAB01 {Rc3ch} 
E1COAXCAB01 n009COAXCAB01 n010COAXCAB01 n007COAXCAB01 n008COAXCAB01 1 
R7COAXCAB01 n010COAXCAB01 RBssCOAXCAB01 {Rc3ch} 
E2COAXCAB01 n008COAXCAB01 LBssCOAXCAB01 n010COAXCAB01 RBssCOAXCAB01 1 
R8COAXCAB01 RBssCOAXCAB01 N050 1e-3 
R9COAXCAB01 LBssCOAXCAB01 N046 1e-3 
* <component=coax_sup>Rs=Rc4h Ls=Lc4h RsG=Rc4g LsG=Lc4g Cp=Cc4sh Rp=Rc4sh k=kc4 Rch=Rc4ch </component>
.param Rs2_COAXCAB02={0.5*Rc4h} Ls2_COAXCAB02={0.5*Lc4h} RsG2_COAXCAB02={0.5*Rc4g} LsG2_COAXCAB02={0.5*Lc4g} 
R1COAXCAB02 N003 n001COAXCAB02 {Rs2_COAXCAB02} 
L1COAXCAB02 n001COAXCAB02 n002COAXCAB02 {Ls2_COAXCAB02} 
L2COAXCAB02 n002COAXCAB02 n003COAXCAB02 {Ls2_COAXCAB02} 
R2COAXCAB02 n003COAXCAB02 n007COAXCAB02 {Rs2_COAXCAB02} 
K1COAXCAB02 L1COAXCAB02 L3COAXCAB02 {kc4} 
R3COAXCAB02 N024 n004COAXCAB02 {RsG2_COAXCAB02} 
L3COAXCAB02 n004COAXCAB02 n005COAXCAB02 {LsG2_COAXCAB02} 
L4COAXCAB02 n005COAXCAB02 n006COAXCAB02 {LsG2_COAXCAB02} 
R4COAXCAB02 n006COAXCAB02 n009COAXCAB02 {RsG2_COAXCAB02} 
K2COAXCAB02 L2COAXCAB02 L4COAXCAB02 {kc4} 
C1COAXCAB02 n002COAXCAB02 n005COAXCAB02 {Cc4sh} 
R5COAXCAB02 n002COAXCAB02 n005COAXCAB02 {Rc4sh} 
R6COAXCAB02 n007COAXCAB02 n008COAXCAB02 {Rc4ch} 
E1COAXCAB02 n009COAXCAB02 n010COAXCAB02 n007COAXCAB02 n008COAXCAB02 1 
R7COAXCAB02 n010COAXCAB02 RBssCOAXCAB02 {Rc4ch} 
E2COAXCAB02 n008COAXCAB02 LBssCOAXCAB02 n010COAXCAB02 RBssCOAXCAB02 1 
R8COAXCAB02 RBssCOAXCAB02 N011 1e-3 
R9COAXCAB02 LBssCOAXCAB02 N004 1e-3 
I1 N003 N024 {Idc} AC {Iac} 0
* <component=coax_Z1>Rs=Rc1h Ls=Lc1h RsG=Rc1g LsG=Lc1g Cp=Cc1sh Rp=Rc1sh k=kc1 Rch=Rc1ch </component>
.param Rs2_COAXCAB03={0.5*Rc1h} Ls2_COAXCAB03={0.5*Lc1h} RsG2_COAXCAB03={0.5*Rc1g} LsG2_COAXCAB03={0.5*Lc1g} 
R1COAXCAB03 N047 n001COAXCAB03 {Rs2_COAXCAB03} 
L1COAXCAB03 n001COAXCAB03 n002COAXCAB03 {Ls2_COAXCAB03} 
L2COAXCAB03 n002COAXCAB03 n003COAXCAB03 {Ls2_COAXCAB03} 
R2COAXCAB03 n003COAXCAB03 n007COAXCAB03 {Rs2_COAXCAB03} 
K1COAXCAB03 L1COAXCAB03 L3COAXCAB03 {kc1} 
R3COAXCAB03 N051 n004COAXCAB03 {RsG2_COAXCAB03} 
L3COAXCAB03 n004COAXCAB03 n005COAXCAB03 {LsG2_COAXCAB03} 
L4COAXCAB03 n005COAXCAB03 n006COAXCAB03 {LsG2_COAXCAB03} 
R4COAXCAB03 n006COAXCAB03 n009COAXCAB03 {RsG2_COAXCAB03} 
K2COAXCAB03 L2COAXCAB03 L4COAXCAB03 {kc1} 
C1COAXCAB03 n002COAXCAB03 n005COAXCAB03 {Cc1sh} 
R5COAXCAB03 n002COAXCAB03 n005COAXCAB03 {Rc1sh} 
R6COAXCAB03 n007COAXCAB03 n008COAXCAB03 {Rc1ch} 
E1COAXCAB03 n009COAXCAB03 n010COAXCAB03 n007COAXCAB03 n008COAXCAB03 1 
R7COAXCAB03 n010COAXCAB03 RBssCOAXCAB03 {Rc1ch} 
E2COAXCAB03 n008COAXCAB03 LBssCOAXCAB03 n010COAXCAB03 RBssCOAXCAB03 1 
R8COAXCAB03 RBssCOAXCAB03 N052 1e-3 
R9COAXCAB03 LBssCOAXCAB03 N048 1e-3 
R1GNDLUG01 N020 n001GNDLUG01 {Rgrd3} 
L1GNDLUG01 n001GNDLUG01 N022 {Lgrd3} 
R1GNDLUG02 N054 n001GNDLUG02 {Rgnd1} 
L1GNDLUG02 n001GNDLUG02 0 {Lgnd1} 
R1GNDLUG03 N037 n001GNDLUG03 {Rsrc} 
L1GNDLUG03 n001GNDLUG03 0 {Lsrc} 
XZ2 N005 N012 N039 N030 N004 N011 N038 N029 NC_01 NC_02 STD4TP3 Rp={Rp2} Lp={Lp2} Rpg={Rp2r} Lpg={Lp2r} kp={kpo2} Cps={Cp2s} Rps={Rp2s} Rc={Rc2} Lc={Lc2} Rcg={Rc2r} Lcg={Lc2r} kc={kco2} Ccs={Cc2s} Rcs={Rc2s} Rs={R2} Ls={L2} Rg={R2g} Lg={L2g} Rb={R2b} Lb={L2b}
R1GNDLUG04 N021 n001GNDLUG04 {Rgnd3} 
L1GNDLUG04 n001GNDLUG04 0 {Lgnd3} 
R1GNDLUG05 N025 n001GNDLUG05 {Rgrd2} 
L1GNDLUG05 n001GNDLUG05 N026 {Lgrd2} 
R1GNDLUG06 N027 n001GNDLUG06 {Rgnd2} 
L1GNDLUG06 n001GNDLUG06 0 {Lgnd2} 
* <component=Hpot_A>Rs=RsHpot_A Ls=LsHpot_A RsG=RsGHpot_A LsG=LsGHpot_A Mlg=MlgHpot_A Cp=CpHpot_A Rp=RpHpot_A RsS=RsSHpot_A LsS=LsSHpot_A Mls=MlsHpot_A Mgs=MgsHpot_A CpS=CpSHpot_A RpS=RpSHpot_A Mll=MllHpot_A Mgg=MggHpot_A Mlg2=Mlg2Hpot_A CpGG=CpGGHpot_A RpGG=RpGGHpot_A </component>
.param Rs2_TWAXSH01={0.5*RsHpot_A} Ls2_TWAXSH01={0.5*LsHpot_A} RsG2_TWAXSH01={0.5*RsGHpot_A} LsG2_TWAXSH01={0.5*LsGHpot_A} RsS2_TWAXSH01={0.5*RsSHpot_A} LsS2_TWAXSH01={0.5*LsSHpot_A} 
.param Rnull_TWAXSH01=1e9 
.param k_lg_TWAXSH01={MlgHpot_A/sqrt(LsHpot_A*LsGHpot_A)} k_ls_TWAXSH01={MlsHpot_A/sqrt(LsHpot_A*LsSHpot_A)} k_gs_TWAXSH01={MgsHpot_A/sqrt(LsGHpot_A*LsSHpot_A)} k_gg_TWAXSH01={MggHpot_A/sqrt(LsGHpot_A*LsGHpot_A)} k_ll_TWAXSH01={MllHpot_A/sqrt(LsHpot_A*LsHpot_A)} k_lg2_TWAXSH01={Mlg2Hpot_A/sqrt(LsHpot_A*LsGHpot_A)} 
L1TWAXSH01 N003TWAXSH01 P001TWAXSH01 {LsG2_TWAXSH01} 
L2TWAXSH01 N004TWAXSH01 P002TWAXSH01 {Ls2_TWAXSH01} 
L3TWAXSH01 P003TWAXSH01 N003TWAXSH01 {LsG2_TWAXSH01} 
L4TWAXSH01 P004TWAXSH01 N004TWAXSH01 {Ls2_TWAXSH01} 
C1TWAXSH01 N003TWAXSH01 N004TWAXSH01 {CpHpot_A} 
R1TWAXSH01 N003TWAXSH01 N004TWAXSH01 {RpHpot_A} 
R2TWAXSH01 P001TWAXSH01 N001 {RsG2_TWAXSH01} 
R3TWAXSH01 P002TWAXSH01 N008 {Rs2_TWAXSH01} 
R4TWAXSH01 N007 P004TWAXSH01 {Rs2_TWAXSH01} 
R5TWAXSH01 NC_04 P003TWAXSH01 {RsG2_TWAXSH01} 
L5TWAXSH01 N001TWAXSH01 P005TWAXSH01 {Ls2_TWAXSH01} 
L6TWAXSH01 N002TWAXSH01 P006TWAXSH01 {LsG2_TWAXSH01} 
L7TWAXSH01 P007TWAXSH01 N001TWAXSH01 {Ls2_TWAXSH01} 
L8TWAXSH01 P008TWAXSH01 N002TWAXSH01 {LsG2_TWAXSH01} 
C2TWAXSH01 N001TWAXSH01 N002TWAXSH01 {CpHpot_A} 
R6TWAXSH01 N001TWAXSH01 N002TWAXSH01 {RpHpot_A} 
R7TWAXSH01 P005TWAXSH01 N015 {Rs2_TWAXSH01} 
R8TWAXSH01 P006TWAXSH01 N019 {RsG2_TWAXSH01} 
R9TWAXSH01 NC_03 P008TWAXSH01 {RsG2_TWAXSH01} 
R10TWAXSH01 N014 P007TWAXSH01 {Rs2_TWAXSH01} 
L9TWAXSH01 CAPTWAXSH01 P009TWAXSH01 {LsS2_TWAXSH01} 
L10TWAXSH01 P010TWAXSH01 CAPTWAXSH01 {LsS2_TWAXSH01} 
R11TWAXSH01 P009TWAXSH01 0 {RsS2_TWAXSH01} 
R12TWAXSH01 NC_05 P010TWAXSH01 {RsS2_TWAXSH01} 
C3TWAXSH01 N002TWAXSH01 CAPTWAXSH01 {CpSHpot_A} 
C4TWAXSH01 CAPTWAXSH01 N003TWAXSH01 {CpSHpot_A} 
R13TWAXSH01 CAPTWAXSH01 N003TWAXSH01 {RpSHpot_A} 
R14TWAXSH01 N002TWAXSH01 CAPTWAXSH01 {RpSHpot_A} 
C5TWAXSH01 N002TWAXSH01 N003TWAXSH01 {CpGGHpot_A} 
R15TWAXSH01 N002TWAXSH01 N003TWAXSH01 {RpGGHpot_A} 
R16TWAXSH01 N015 N019 {Rnull_TWAXSH01} 
R17TWAXSH01 N019 0 {Rnull_TWAXSH01} 
R18TWAXSH01 0 N001 {Rnull_TWAXSH01} 
R19TWAXSH01 N001 N008 {Rnull_TWAXSH01} 
R20TWAXSH01 NC_04 N007 {Rnull_TWAXSH01} 
R21TWAXSH01 NC_05 NC_04 {Rnull_TWAXSH01} 
R22TWAXSH01 NC_03 NC_05 {Rnull_TWAXSH01} 
R23TWAXSH01 N014 NC_03 {Rnull_TWAXSH01} 
KlaTWAXSH01 L5TWAXSH01 L6TWAXSH01 {k_lg_TWAXSH01} 
KraTWAXSH01 L7TWAXSH01 L8TWAXSH01 {k_lg_TWAXSH01} 
KlbTWAXSH01 L1TWAXSH01 L2TWAXSH01 {k_lg_TWAXSH01} 
KrbTWAXSH01 L3TWAXSH01 L4TWAXSH01 {k_lg_TWAXSH01} 
KllsaTWAXSH01 L5TWAXSH01 L9TWAXSH01 {k_ls_TWAXSH01} 
KlgsaTWAXSH01 L6TWAXSH01 L9TWAXSH01 {k_gs_TWAXSH01} 
KlgsbTWAXSH01 L1TWAXSH01 L9TWAXSH01 {k_gs_TWAXSH01} 
KllsbTWAXSH01 L2TWAXSH01 L9TWAXSH01 {k_ls_TWAXSH01} 
KlggTWAXSH01 L6TWAXSH01 L1TWAXSH01 {k_gg_TWAXSH01} 
KlllTWAXSH01 L5TWAXSH01 L2TWAXSH01 {k_ll_TWAXSH01} 
KlglTWAXSH01 L6TWAXSH01 L2TWAXSH01 {k_lg2_TWAXSH01} 
Klgl2TWAXSH01 L5TWAXSH01 L1TWAXSH01 {k_lg2_TWAXSH01} 
KrlsaTWAXSH01 L7TWAXSH01 L10TWAXSH01 {k_ls_TWAXSH01} 
KrgsaTWAXSH01 L8TWAXSH01 L10TWAXSH01 {k_gs_TWAXSH01} 
KrgsbTWAXSH01 L3TWAXSH01 L10TWAXSH01 {k_gs_TWAXSH01} 
KrlsbTWAXSH01 L4TWAXSH01 L10TWAXSH01 {k_ls_TWAXSH01} 
KrggTWAXSH01 L8TWAXSH01 L3TWAXSH01 {k_gg_TWAXSH01} 
KrllTWAXSH01 L7TWAXSH01 L4TWAXSH01 {k_ll_TWAXSH01} 
KrglTWAXSH01 L8TWAXSH01 L4TWAXSH01 {k_lg2_TWAXSH01} 
Krgl2TWAXSH01 L7TWAXSH01 L3TWAXSH01 {k_lg2_TWAXSH01} 
* <component=Lpot_A>Rs=RsLpot_A Ls=LsLpot_A RsG=RsGLpot_A LsG=LsGLpot_A Mlg=MlgLpot_A Cp=CpLpot_A Rp=RpLpot_A RsS=RsSLpot_A LsS=LsSLpot_A Mls=MlsLpot_A Mgs=MgsLpot_A CpS=CpSLpot_A RpS=RpSLpot_A Mll=MllLpot_A Mgg=MggLpot_A Mlg2=Mlg2Lpot_A CpGG=CpGGLpot_A RpGG=RpGGLpot_A </component>
.param Rs2_TWAXSH02={0.5*RsLpot_A} Ls2_TWAXSH02={0.5*LsLpot_A} RsG2_TWAXSH02={0.5*RsGLpot_A} LsG2_TWAXSH02={0.5*LsGLpot_A} RsS2_TWAXSH02={0.5*RsSLpot_A} LsS2_TWAXSH02={0.5*LsSLpot_A} 
.param Rnull_TWAXSH02=1e9 
.param k_lg_TWAXSH02={MlgLpot_A/sqrt(LsLpot_A*LsGLpot_A)} k_ls_TWAXSH02={MlsLpot_A/sqrt(LsLpot_A*LsSLpot_A)} k_gs_TWAXSH02={MgsLpot_A/sqrt(LsGLpot_A*LsSLpot_A)} k_gg_TWAXSH02={MggLpot_A/sqrt(LsGLpot_A*LsGLpot_A)} k_ll_TWAXSH02={MllLpot_A/sqrt(LsLpot_A*LsLpot_A)} k_lg2_TWAXSH02={Mlg2Lpot_A/sqrt(LsLpot_A*LsGLpot_A)} 
L1TWAXSH02 N003TWAXSH02 P001TWAXSH02 {LsG2_TWAXSH02} 
L2TWAXSH02 N004TWAXSH02 P002TWAXSH02 {Ls2_TWAXSH02} 
L3TWAXSH02 P003TWAXSH02 N003TWAXSH02 {LsG2_TWAXSH02} 
L4TWAXSH02 P004TWAXSH02 N004TWAXSH02 {Ls2_TWAXSH02} 
C1TWAXSH02 N003TWAXSH02 N004TWAXSH02 {CpLpot_A} 
R1TWAXSH02 N003TWAXSH02 N004TWAXSH02 {RpLpot_A} 
R2TWAXSH02 P001TWAXSH02 NC_07 {RsG2_TWAXSH02} 
R3TWAXSH02 P002TWAXSH02 N040 {Rs2_TWAXSH02} 
R4TWAXSH02 N041 P004TWAXSH02 {Rs2_TWAXSH02} 
R5TWAXSH02 N044 P003TWAXSH02 {RsG2_TWAXSH02} 
L5TWAXSH02 N001TWAXSH02 P005TWAXSH02 {Ls2_TWAXSH02} 
L6TWAXSH02 N002TWAXSH02 P006TWAXSH02 {LsG2_TWAXSH02} 
L7TWAXSH02 P007TWAXSH02 N001TWAXSH02 {Ls2_TWAXSH02} 
L8TWAXSH02 P008TWAXSH02 N002TWAXSH02 {LsG2_TWAXSH02} 
C2TWAXSH02 N001TWAXSH02 N002TWAXSH02 {CpLpot_A} 
R6TWAXSH02 N001TWAXSH02 N002TWAXSH02 {RpLpot_A} 
R7TWAXSH02 P005TWAXSH02 N032 {Rs2_TWAXSH02} 
R8TWAXSH02 P006TWAXSH02 NC_06 {RsG2_TWAXSH02} 
R9TWAXSH02 N028 P008TWAXSH02 {RsG2_TWAXSH02} 
R10TWAXSH02 N033 P007TWAXSH02 {Rs2_TWAXSH02} 
L9TWAXSH02 CAPTWAXSH02 P009TWAXSH02 {LsS2_TWAXSH02} 
L10TWAXSH02 P010TWAXSH02 CAPTWAXSH02 {LsS2_TWAXSH02} 
R11TWAXSH02 P009TWAXSH02 NC_08 {RsS2_TWAXSH02} 
R12TWAXSH02 0 P010TWAXSH02 {RsS2_TWAXSH02} 
C3TWAXSH02 N002TWAXSH02 CAPTWAXSH02 {CpSLpot_A} 
C4TWAXSH02 CAPTWAXSH02 N003TWAXSH02 {CpSLpot_A} 
R13TWAXSH02 CAPTWAXSH02 N003TWAXSH02 {RpSLpot_A} 
R14TWAXSH02 N002TWAXSH02 CAPTWAXSH02 {RpSLpot_A} 
C5TWAXSH02 N002TWAXSH02 N003TWAXSH02 {CpGGLpot_A} 
R15TWAXSH02 N002TWAXSH02 N003TWAXSH02 {RpGGLpot_A} 
R16TWAXSH02 N032 NC_06 {Rnull_TWAXSH02} 
R17TWAXSH02 NC_06 NC_08 {Rnull_TWAXSH02} 
R18TWAXSH02 NC_08 NC_07 {Rnull_TWAXSH02} 
R19TWAXSH02 NC_07 N040 {Rnull_TWAXSH02} 
R20TWAXSH02 N044 N041 {Rnull_TWAXSH02} 
R21TWAXSH02 0 N044 {Rnull_TWAXSH02} 
R22TWAXSH02 N028 0 {Rnull_TWAXSH02} 
R23TWAXSH02 N033 N028 {Rnull_TWAXSH02} 
KlaTWAXSH02 L5TWAXSH02 L6TWAXSH02 {k_lg_TWAXSH02} 
KraTWAXSH02 L7TWAXSH02 L8TWAXSH02 {k_lg_TWAXSH02} 
KlbTWAXSH02 L1TWAXSH02 L2TWAXSH02 {k_lg_TWAXSH02} 
KrbTWAXSH02 L3TWAXSH02 L4TWAXSH02 {k_lg_TWAXSH02} 
KllsaTWAXSH02 L5TWAXSH02 L9TWAXSH02 {k_ls_TWAXSH02} 
KlgsaTWAXSH02 L6TWAXSH02 L9TWAXSH02 {k_gs_TWAXSH02} 
KlgsbTWAXSH02 L1TWAXSH02 L9TWAXSH02 {k_gs_TWAXSH02} 
KllsbTWAXSH02 L2TWAXSH02 L9TWAXSH02 {k_ls_TWAXSH02} 
KlggTWAXSH02 L6TWAXSH02 L1TWAXSH02 {k_gg_TWAXSH02} 
KlllTWAXSH02 L5TWAXSH02 L2TWAXSH02 {k_ll_TWAXSH02} 
KlglTWAXSH02 L6TWAXSH02 L2TWAXSH02 {k_lg2_TWAXSH02} 
Klgl2TWAXSH02 L5TWAXSH02 L1TWAXSH02 {k_lg2_TWAXSH02} 
KrlsaTWAXSH02 L7TWAXSH02 L10TWAXSH02 {k_ls_TWAXSH02} 
KrgsaTWAXSH02 L8TWAXSH02 L10TWAXSH02 {k_gs_TWAXSH02} 
KrgsbTWAXSH02 L3TWAXSH02 L10TWAXSH02 {k_gs_TWAXSH02} 
KrlsbTWAXSH02 L4TWAXSH02 L10TWAXSH02 {k_ls_TWAXSH02} 
KrggTWAXSH02 L8TWAXSH02 L3TWAXSH02 {k_gg_TWAXSH02} 
KrllTWAXSH02 L7TWAXSH02 L4TWAXSH02 {k_ll_TWAXSH02} 
KrglTWAXSH02 L8TWAXSH02 L4TWAXSH02 {k_lg2_TWAXSH02} 
Krgl2TWAXSH02 L7TWAXSH02 L3TWAXSH02 {k_lg2_TWAXSH02} 
* <component=buf_hpot>CgA=CgA_buf_hpot RgA=RgA_buf_hpot CgB=CgB_buf_hpot RgB=RgB_buf_hpot LoA=LoA_buf_hpot RoA=RoA_buf_hpot LoB=LoB_buf_hpot RoB=RoB_buf_hpot </component>
Xbuf_hpot N008 N001 N015 N019 N009 N002 N016 N020 0 DUAL_EPBUF CgA={CgA_buf_hpot} RgA={RgA_buf_hpot} CgB={CgB_buf_hpot} RgB={RgB_buf_hpot} LoA={LoA_buf_hpot} RoA={RoA_buf_hpot} LoB={LoB_buf_hpot} RoB={RoB_buf_hpot} 
* <component=buf_lpot>CgA=CgA_buf_lpot RgA=RgA_buf_lpot CgB=CgB_buf_lpot RgB=RgB_buf_lpot LoA=LoA_buf_lpot RoA=RoA_buf_lpot LoB=LoB_buf_lpot RoB=RoB_buf_lpot </component>
Xbuf_lpot N042 N045 N034 N025 N041 N044 N033 N028 0 DUAL_EPBUF CgA={CgA_buf_lpot} RgA={RgA_buf_lpot} CgB={CgB_buf_lpot} RgB={RgB_buf_lpot} LoA={LoA_buf_lpot} RoA={RoA_buf_lpot} LoB={LoB_buf_lpot} RoB={RoB_buf_lpot} 
* <component=Hpot_B>Rs=RsHpot_B Ls=LsHpot_B RsG=RsGHpot_B LsG=LsGHpot_B Mlg=MlgHpot_B Cp=CpHpot_B Rp=RpHpot_B RsS=RsSHpot_B LsS=LsSHpot_B Mls=MlsHpot_B Mgs=MgsHpot_B CpS=CpSHpot_B RpS=RpSHpot_B Mll=MllHpot_B Mgg=MggHpot_B Mlg2=Mlg2Hpot_B CpGG=CpGGHpot_B RpGG=RpGGHpot_B </component>
.param Rs2_TWAXSH03={0.5*RsHpot_B} Ls2_TWAXSH03={0.5*LsHpot_B} RsG2_TWAXSH03={0.5*RsGHpot_B} LsG2_TWAXSH03={0.5*LsGHpot_B} RsS2_TWAXSH03={0.5*RsSHpot_B} LsS2_TWAXSH03={0.5*LsSHpot_B} 
.param Rnull_TWAXSH03=1e9 
.param k_lg_TWAXSH03={MlgHpot_B/sqrt(LsHpot_B*LsGHpot_B)} k_ls_TWAXSH03={MlsHpot_B/sqrt(LsHpot_B*LsSHpot_B)} k_gs_TWAXSH03={MgsHpot_B/sqrt(LsGHpot_B*LsSHpot_B)} k_gg_TWAXSH03={MggHpot_B/sqrt(LsGHpot_B*LsGHpot_B)} k_ll_TWAXSH03={MllHpot_B/sqrt(LsHpot_B*LsHpot_B)} k_lg2_TWAXSH03={Mlg2Hpot_B/sqrt(LsHpot_B*LsGHpot_B)} 
L1TWAXSH03 N003TWAXSH03 P001TWAXSH03 {LsG2_TWAXSH03} 
L2TWAXSH03 N004TWAXSH03 P002TWAXSH03 {Ls2_TWAXSH03} 
L3TWAXSH03 P003TWAXSH03 N003TWAXSH03 {LsG2_TWAXSH03} 
L4TWAXSH03 P004TWAXSH03 N004TWAXSH03 {Ls2_TWAXSH03} 
C1TWAXSH03 N003TWAXSH03 N004TWAXSH03 {CpHpot_B} 
R1TWAXSH03 N003TWAXSH03 N004TWAXSH03 {RpHpot_B} 
R2TWAXSH03 P001TWAXSH03 NC_10 {RsG2_TWAXSH03} 
R3TWAXSH03 P002TWAXSH03 U3 {Rs2_TWAXSH03} 
R4TWAXSH03 N009 P004TWAXSH03 {Rs2_TWAXSH03} 
R5TWAXSH03 N002 P003TWAXSH03 {RsG2_TWAXSH03} 
L5TWAXSH03 N001TWAXSH03 P005TWAXSH03 {Ls2_TWAXSH03} 
L6TWAXSH03 N002TWAXSH03 P006TWAXSH03 {LsG2_TWAXSH03} 
L7TWAXSH03 P007TWAXSH03 N001TWAXSH03 {Ls2_TWAXSH03} 
L8TWAXSH03 P008TWAXSH03 N002TWAXSH03 {LsG2_TWAXSH03} 
C2TWAXSH03 N001TWAXSH03 N002TWAXSH03 {CpHpot_B} 
R6TWAXSH03 N001TWAXSH03 N002TWAXSH03 {RpHpot_B} 
R7TWAXSH03 P005TWAXSH03 N017 {Rs2_TWAXSH03} 
R8TWAXSH03 P006TWAXSH03 NC_09 {RsG2_TWAXSH03} 
R9TWAXSH03 N020 P008TWAXSH03 {RsG2_TWAXSH03} 
R10TWAXSH03 N016 P007TWAXSH03 {Rs2_TWAXSH03} 
L9TWAXSH03 CAPTWAXSH03 P009TWAXSH03 {LsS2_TWAXSH03} 
L10TWAXSH03 P010TWAXSH03 CAPTWAXSH03 {LsS2_TWAXSH03} 
R11TWAXSH03 P009TWAXSH03 NC_11 {RsS2_TWAXSH03} 
R12TWAXSH03 0 P010TWAXSH03 {RsS2_TWAXSH03} 
C3TWAXSH03 N002TWAXSH03 CAPTWAXSH03 {CpSHpot_B} 
C4TWAXSH03 CAPTWAXSH03 N003TWAXSH03 {CpSHpot_B} 
R13TWAXSH03 CAPTWAXSH03 N003TWAXSH03 {RpSHpot_B} 
R14TWAXSH03 N002TWAXSH03 CAPTWAXSH03 {RpSHpot_B} 
C5TWAXSH03 N002TWAXSH03 N003TWAXSH03 {CpGGHpot_B} 
R15TWAXSH03 N002TWAXSH03 N003TWAXSH03 {RpGGHpot_B} 
R16TWAXSH03 N017 NC_09 {Rnull_TWAXSH03} 
R17TWAXSH03 NC_09 NC_11 {Rnull_TWAXSH03} 
R18TWAXSH03 NC_11 NC_10 {Rnull_TWAXSH03} 
R19TWAXSH03 NC_10 U3 {Rnull_TWAXSH03} 
R20TWAXSH03 N002 N009 {Rnull_TWAXSH03} 
R21TWAXSH03 0 N002 {Rnull_TWAXSH03} 
R22TWAXSH03 N020 0 {Rnull_TWAXSH03} 
R23TWAXSH03 N016 N020 {Rnull_TWAXSH03} 
KlaTWAXSH03 L5TWAXSH03 L6TWAXSH03 {k_lg_TWAXSH03} 
KraTWAXSH03 L7TWAXSH03 L8TWAXSH03 {k_lg_TWAXSH03} 
KlbTWAXSH03 L1TWAXSH03 L2TWAXSH03 {k_lg_TWAXSH03} 
KrbTWAXSH03 L3TWAXSH03 L4TWAXSH03 {k_lg_TWAXSH03} 
KllsaTWAXSH03 L5TWAXSH03 L9TWAXSH03 {k_ls_TWAXSH03} 
KlgsaTWAXSH03 L6TWAXSH03 L9TWAXSH03 {k_gs_TWAXSH03} 
KlgsbTWAXSH03 L1TWAXSH03 L9TWAXSH03 {k_gs_TWAXSH03} 
KllsbTWAXSH03 L2TWAXSH03 L9TWAXSH03 {k_ls_TWAXSH03} 
KlggTWAXSH03 L6TWAXSH03 L1TWAXSH03 {k_gg_TWAXSH03} 
KlllTWAXSH03 L5TWAXSH03 L2TWAXSH03 {k_ll_TWAXSH03} 
KlglTWAXSH03 L6TWAXSH03 L2TWAXSH03 {k_lg2_TWAXSH03} 
Klgl2TWAXSH03 L5TWAXSH03 L1TWAXSH03 {k_lg2_TWAXSH03} 
KrlsaTWAXSH03 L7TWAXSH03 L10TWAXSH03 {k_ls_TWAXSH03} 
KrgsaTWAXSH03 L8TWAXSH03 L10TWAXSH03 {k_gs_TWAXSH03} 
KrgsbTWAXSH03 L3TWAXSH03 L10TWAXSH03 {k_gs_TWAXSH03} 
KrlsbTWAXSH03 L4TWAXSH03 L10TWAXSH03 {k_ls_TWAXSH03} 
KrggTWAXSH03 L8TWAXSH03 L3TWAXSH03 {k_gg_TWAXSH03} 
KrllTWAXSH03 L7TWAXSH03 L4TWAXSH03 {k_ll_TWAXSH03} 
KrglTWAXSH03 L8TWAXSH03 L4TWAXSH03 {k_lg2_TWAXSH03} 
Krgl2TWAXSH03 L7TWAXSH03 L3TWAXSH03 {k_lg2_TWAXSH03} 
* <component=Lpot_B>Rs=RsLpot_B Ls=LsLpot_B RsG=RsGLpot_B LsG=LsGLpot_B Mlg=MlgLpot_B Cp=CpLpot_B Rp=RpLpot_B RsS=RsSLpot_B LsS=LsSLpot_B Mls=MlsLpot_B Mgs=MgsLpot_B CpS=CpSLpot_B RpS=RpSLpot_B Mll=MllLpot_B Mgg=MggLpot_B Mlg2=Mlg2Lpot_B CpGG=CpGGLpot_B RpGG=RpGGLpot_B </component>
.param Rs2_TWAXSH04={0.5*RsLpot_B} Ls2_TWAXSH04={0.5*LsLpot_B} RsG2_TWAXSH04={0.5*RsGLpot_B} LsG2_TWAXSH04={0.5*LsGLpot_B} RsS2_TWAXSH04={0.5*RsSLpot_B} LsS2_TWAXSH04={0.5*LsSLpot_B} 
.param Rnull_TWAXSH04=1e9 
.param k_lg_TWAXSH04={MlgLpot_B/sqrt(LsLpot_B*LsGLpot_B)} k_ls_TWAXSH04={MlsLpot_B/sqrt(LsLpot_B*LsSLpot_B)} k_gs_TWAXSH04={MgsLpot_B/sqrt(LsGLpot_B*LsSLpot_B)} k_gg_TWAXSH04={MggLpot_B/sqrt(LsGLpot_B*LsGLpot_B)} k_ll_TWAXSH04={MllLpot_B/sqrt(LsLpot_B*LsLpot_B)} k_lg2_TWAXSH04={Mlg2Lpot_B/sqrt(LsLpot_B*LsGLpot_B)} 
L1TWAXSH04 N003TWAXSH04 P001TWAXSH04 {LsG2_TWAXSH04} 
L2TWAXSH04 N004TWAXSH04 P002TWAXSH04 {Ls2_TWAXSH04} 
L3TWAXSH04 P003TWAXSH04 N003TWAXSH04 {LsG2_TWAXSH04} 
L4TWAXSH04 P004TWAXSH04 N004TWAXSH04 {Ls2_TWAXSH04} 
C1TWAXSH04 N003TWAXSH04 N004TWAXSH04 {CpLpot_B} 
R1TWAXSH04 N003TWAXSH04 N004TWAXSH04 {RpLpot_B} 
R2TWAXSH04 P001TWAXSH04 N045 {RsG2_TWAXSH04} 
R3TWAXSH04 P002TWAXSH04 N042 {Rs2_TWAXSH04} 
R4TWAXSH04 U2 P004TWAXSH04 {Rs2_TWAXSH04} 
R5TWAXSH04 NC_13 P003TWAXSH04 {RsG2_TWAXSH04} 
L5TWAXSH04 N001TWAXSH04 P005TWAXSH04 {Ls2_TWAXSH04} 
L6TWAXSH04 N002TWAXSH04 P006TWAXSH04 {LsG2_TWAXSH04} 
L7TWAXSH04 P007TWAXSH04 N001TWAXSH04 {Ls2_TWAXSH04} 
L8TWAXSH04 P008TWAXSH04 N002TWAXSH04 {LsG2_TWAXSH04} 
C2TWAXSH04 N001TWAXSH04 N002TWAXSH04 {CpLpot_B} 
R6TWAXSH04 N001TWAXSH04 N002TWAXSH04 {RpLpot_B} 
R7TWAXSH04 P005TWAXSH04 N034 {Rs2_TWAXSH04} 
R8TWAXSH04 P006TWAXSH04 N025 {RsG2_TWAXSH04} 
R9TWAXSH04 NC_12 P008TWAXSH04 {RsG2_TWAXSH04} 
R10TWAXSH04 N035 P007TWAXSH04 {Rs2_TWAXSH04} 
L9TWAXSH04 CAPTWAXSH04 P009TWAXSH04 {LsS2_TWAXSH04} 
L10TWAXSH04 P010TWAXSH04 CAPTWAXSH04 {LsS2_TWAXSH04} 
R11TWAXSH04 P009TWAXSH04 0 {RsS2_TWAXSH04} 
R12TWAXSH04 NC_14 P010TWAXSH04 {RsS2_TWAXSH04} 
C3TWAXSH04 N002TWAXSH04 CAPTWAXSH04 {CpSLpot_B} 
C4TWAXSH04 CAPTWAXSH04 N003TWAXSH04 {CpSLpot_B} 
R13TWAXSH04 CAPTWAXSH04 N003TWAXSH04 {RpSLpot_B} 
R14TWAXSH04 N002TWAXSH04 CAPTWAXSH04 {RpSLpot_B} 
C5TWAXSH04 N002TWAXSH04 N003TWAXSH04 {CpGGLpot_B} 
R15TWAXSH04 N002TWAXSH04 N003TWAXSH04 {RpGGLpot_B} 
R16TWAXSH04 N034 N025 {Rnull_TWAXSH04} 
R17TWAXSH04 N025 0 {Rnull_TWAXSH04} 
R18TWAXSH04 0 N045 {Rnull_TWAXSH04} 
R19TWAXSH04 N045 N042 {Rnull_TWAXSH04} 
R20TWAXSH04 NC_13 U2 {Rnull_TWAXSH04} 
R21TWAXSH04 NC_14 NC_13 {Rnull_TWAXSH04} 
R22TWAXSH04 NC_12 NC_14 {Rnull_TWAXSH04} 
R23TWAXSH04 N035 NC_12 {Rnull_TWAXSH04} 
KlaTWAXSH04 L5TWAXSH04 L6TWAXSH04 {k_lg_TWAXSH04} 
KraTWAXSH04 L7TWAXSH04 L8TWAXSH04 {k_lg_TWAXSH04} 
KlbTWAXSH04 L1TWAXSH04 L2TWAXSH04 {k_lg_TWAXSH04} 
KrbTWAXSH04 L3TWAXSH04 L4TWAXSH04 {k_lg_TWAXSH04} 
KllsaTWAXSH04 L5TWAXSH04 L9TWAXSH04 {k_ls_TWAXSH04} 
KlgsaTWAXSH04 L6TWAXSH04 L9TWAXSH04 {k_gs_TWAXSH04} 
KlgsbTWAXSH04 L1TWAXSH04 L9TWAXSH04 {k_gs_TWAXSH04} 
KllsbTWAXSH04 L2TWAXSH04 L9TWAXSH04 {k_ls_TWAXSH04} 
KlggTWAXSH04 L6TWAXSH04 L1TWAXSH04 {k_gg_TWAXSH04} 
KlllTWAXSH04 L5TWAXSH04 L2TWAXSH04 {k_ll_TWAXSH04} 
KlglTWAXSH04 L6TWAXSH04 L2TWAXSH04 {k_lg2_TWAXSH04} 
Klgl2TWAXSH04 L5TWAXSH04 L1TWAXSH04 {k_lg2_TWAXSH04} 
KrlsaTWAXSH04 L7TWAXSH04 L10TWAXSH04 {k_ls_TWAXSH04} 
KrgsaTWAXSH04 L8TWAXSH04 L10TWAXSH04 {k_gs_TWAXSH04} 
KrgsbTWAXSH04 L3TWAXSH04 L10TWAXSH04 {k_gs_TWAXSH04} 
KrlsbTWAXSH04 L4TWAXSH04 L10TWAXSH04 {k_ls_TWAXSH04} 
KrggTWAXSH04 L8TWAXSH04 L3TWAXSH04 {k_gg_TWAXSH04} 
KrllTWAXSH04 L7TWAXSH04 L4TWAXSH04 {k_ll_TWAXSH04} 
KrglTWAXSH04 L8TWAXSH04 L4TWAXSH04 {k_lg2_TWAXSH04} 
Krgl2TWAXSH04 L7TWAXSH04 L3TWAXSH04 {k_lg2_TWAXSH04} 
* <component=ADC3>Ci=Ca3in Ri=Ra3in Clg=Ca3lg Rlg=Ra3lg Cgs=Ca3gs Rgs=Ra3gs guard=grda3 </component>
XADC3 N010 N018 N022 N021 U3_adc_high U3_adc_low DIG3458 Ci={Ca3in} Ri={Ra3in} Clg={Ca3lg} Rlg={Ra3lg} Cgs={Ca3gs} Rgs={Ra3gs} guard={grda3}  
* <component=ADC2>Ci=Ca2in Ri=Ra2in Clg=Ca2lg Rlg=Ra2lg Cgs=Ca2gs Rgs=Ra2gs guard=grda2 </component>
XADC2 N043 N036 N026 N027 U2_adc_high U2_adc_low DIG3458 Ci={Ca2in} Ri={Ra2in} Clg={Ca2lg} Rlg={Ra2lg} Cgs={Ca2gs} Rgs={Ra2gs} guard={grda2}  
* <component=ADC1>Ci=Ca1in Ri=Ra1in Clg=Ca1lg Rlg=Ra1lg Cgs=Ca1gs Rgs=Ra1gs guard=grda1 </component>
XADC1 N049 N053 N055 N054 U1_adc_high U1_adc_low DIG3458 Ci={Ca1in} Ri={Ra1in} Clg={Ca1lg} Rlg={Ra1lg} Cgs={Ca1gs} Rgs={Ra1gs} guard={grda1}  
R1GNDLUG07 N050 n001GNDLUG07 {Rgrd2} 
L1GNDLUG07 n001GNDLUG07 N055 {Lgrd2} 
C1 N024 N037 {Cpsrc}
R1 N024 N037 {Rpsrc}
R1GNDLUG08 N050 n001GNDLUG08 {Rgref} 
L1GNDLUG08 n001GNDLUG08 0 {Lgref} 
* <component=wa3hi>Ls=Rwa3hi Rs=Lwa3hi </component>
R1GNDLUG09 U3 n001GNDLUG09 {Lwa3hi} 
L1GNDLUG09 n001GNDLUG09 N010 {Rwa3hi} 
* <component=wa3lo>Ls=Rwa3lo Rs=Lwa3lo </component>
R1GNDLUG10 N017 n001GNDLUG10 {Lwa3lo} 
L1GNDLUG10 n001GNDLUG10 N018 {Rwa3lo} 
* <component=wa2hi>Ls=Rwa2hi Rs=Lwa2hi </component>
R1GNDLUG11 U2 n001GNDLUG11 {Lwa2hi} 
L1GNDLUG11 n001GNDLUG11 N043 {Rwa2hi} 
* <component=wa2lo>Ls=Rwa2lo Rs=Lwa2lo </component>
R1GNDLUG12 N035 n001GNDLUG12 {Lwa2lo} 
L1GNDLUG12 n001GNDLUG12 N036 {Rwa2lo} 
* <component=wa1hi>Ls=Rwa1hi Rs=Lwa1hi </component>
R1GNDLUG13 N048 n001GNDLUG13 {Lwa1hi} 
L1GNDLUG13 n001GNDLUG13 N049 {Rwa1hi} 
* <component=wa1lo>Ls=Rwa1lo Rs=Lwa1lo </component>
R1GNDLUG14 N052 n001GNDLUG14 {Lwa1lo} 
L1GNDLUG14 n001GNDLUG14 N053 {Rwa1lo} 
* <component=coax_2hi>Rs=Rccoax_2hih Ls=Lccoax_2hih RsG=Rccoax_2hig LsG=Lccoax_2hig Cp=Cccoax_2hish Rp=Rccoax_2hish k=kccoax_2hi Rch=Rccoax_2hich </component>
.param Rs2_COAXCAB04={0.5*Rccoax_2hih} Ls2_COAXCAB04={0.5*Lccoax_2hih} RsG2_COAXCAB04={0.5*Rccoax_2hig} LsG2_COAXCAB04={0.5*Lccoax_2hig} 
R1COAXCAB04 N005 n001COAXCAB04 {Rs2_COAXCAB04} 
L1COAXCAB04 n001COAXCAB04 n002COAXCAB04 {Ls2_COAXCAB04} 
L2COAXCAB04 n002COAXCAB04 n003COAXCAB04 {Ls2_COAXCAB04} 
R2COAXCAB04 n003COAXCAB04 n007COAXCAB04 {Rs2_COAXCAB04} 
K1COAXCAB04 L1COAXCAB04 L3COAXCAB04 {kccoax_2hi} 
R3COAXCAB04 N012 n004COAXCAB04 {RsG2_COAXCAB04} 
L3COAXCAB04 n004COAXCAB04 n005COAXCAB04 {LsG2_COAXCAB04} 
L4COAXCAB04 n005COAXCAB04 n006COAXCAB04 {LsG2_COAXCAB04} 
R4COAXCAB04 n006COAXCAB04 n009COAXCAB04 {RsG2_COAXCAB04} 
K2COAXCAB04 L2COAXCAB04 L4COAXCAB04 {kccoax_2hi} 
C1COAXCAB04 n002COAXCAB04 n005COAXCAB04 {Cccoax_2hish} 
R5COAXCAB04 n002COAXCAB04 n005COAXCAB04 {Rccoax_2hish} 
R6COAXCAB04 n007COAXCAB04 n008COAXCAB04 {Rccoax_2hich} 
E1COAXCAB04 n009COAXCAB04 n010COAXCAB04 n007COAXCAB04 n008COAXCAB04 1 
R7COAXCAB04 n010COAXCAB04 RBssCOAXCAB04 {Rccoax_2hich} 
E2COAXCAB04 n008COAXCAB04 LBssCOAXCAB04 n010COAXCAB04 RBssCOAXCAB04 1 
R8COAXCAB04 RBssCOAXCAB04 N013 1e-3 
R9COAXCAB04 LBssCOAXCAB04 N006 1e-3 
* <component=coax_2lo>Rs=Rccoax_2loh Ls=Lccoax_2loh RsG=Rccoax_2log LsG=Lccoax_2log Cp=Cccoax_2losh Rp=Rccoax_2losh k=kccoax_2lo Rch=Rccoax_2loch </component>
.param Rs2_COAXCAB05={0.5*Rccoax_2loh} Ls2_COAXCAB05={0.5*Lccoax_2loh} RsG2_COAXCAB05={0.5*Rccoax_2log} LsG2_COAXCAB05={0.5*Lccoax_2log} 
R1COAXCAB05 N039 n001COAXCAB05 {Rs2_COAXCAB05} 
L1COAXCAB05 n001COAXCAB05 n002COAXCAB05 {Ls2_COAXCAB05} 
L2COAXCAB05 n002COAXCAB05 n003COAXCAB05 {Ls2_COAXCAB05} 
R2COAXCAB05 n003COAXCAB05 n007COAXCAB05 {Rs2_COAXCAB05} 
K1COAXCAB05 L1COAXCAB05 L3COAXCAB05 {kccoax_2lo} 
R3COAXCAB05 N030 n004COAXCAB05 {RsG2_COAXCAB05} 
L3COAXCAB05 n004COAXCAB05 n005COAXCAB05 {LsG2_COAXCAB05} 
L4COAXCAB05 n005COAXCAB05 n006COAXCAB05 {LsG2_COAXCAB05} 
R4COAXCAB05 n006COAXCAB05 n009COAXCAB05 {RsG2_COAXCAB05} 
K2COAXCAB05 L2COAXCAB05 L4COAXCAB05 {kccoax_2lo} 
C1COAXCAB05 n002COAXCAB05 n005COAXCAB05 {Cccoax_2losh} 
R5COAXCAB05 n002COAXCAB05 n005COAXCAB05 {Rccoax_2losh} 
R6COAXCAB05 n007COAXCAB05 n008COAXCAB05 {Rccoax_2loch} 
E1COAXCAB05 n009COAXCAB05 n010COAXCAB05 n007COAXCAB05 n008COAXCAB05 1 
R7COAXCAB05 n010COAXCAB05 RBssCOAXCAB05 {Rccoax_2loch} 
E2COAXCAB05 n008COAXCAB05 LBssCOAXCAB05 n010COAXCAB05 RBssCOAXCAB05 1 
R8COAXCAB05 RBssCOAXCAB05 N031 1e-3 
R9COAXCAB05 LBssCOAXCAB05 N023 1e-3 
* <component=coax_2live>Rs=Rccoax_2liveh Ls=Lccoax_2liveh RsG=Rccoax_2liveg LsG=Lccoax_2liveg Cp=Cccoax_2livesh Rp=Rccoax_2livesh k=kccoax_2live Rch=Rccoax_2livech </component>
.param Rs2_COAXCAB06={0.5*Rccoax_2liveh} Ls2_COAXCAB06={0.5*Lccoax_2liveh} RsG2_COAXCAB06={0.5*Rccoax_2liveg} LsG2_COAXCAB06={0.5*Lccoax_2liveg} 
R1COAXCAB06 N006 n001COAXCAB06 {Rs2_COAXCAB06} 
L1COAXCAB06 n001COAXCAB06 n002COAXCAB06 {Ls2_COAXCAB06} 
L2COAXCAB06 n002COAXCAB06 n003COAXCAB06 {Ls2_COAXCAB06} 
R2COAXCAB06 n003COAXCAB06 n007COAXCAB06 {Rs2_COAXCAB06} 
K1COAXCAB06 L1COAXCAB06 L3COAXCAB06 {kccoax_2live} 
R3COAXCAB06 N023 n004COAXCAB06 {RsG2_COAXCAB06} 
L3COAXCAB06 n004COAXCAB06 n005COAXCAB06 {LsG2_COAXCAB06} 
L4COAXCAB06 n005COAXCAB06 n006COAXCAB06 {LsG2_COAXCAB06} 
R4COAXCAB06 n006COAXCAB06 n009COAXCAB06 {RsG2_COAXCAB06} 
K2COAXCAB06 L2COAXCAB06 L4COAXCAB06 {kccoax_2live} 
C1COAXCAB06 n002COAXCAB06 n005COAXCAB06 {Cccoax_2livesh} 
R5COAXCAB06 n002COAXCAB06 n005COAXCAB06 {Rccoax_2livesh} 
R6COAXCAB06 n007COAXCAB06 n008COAXCAB06 {Rccoax_2livech} 
E1COAXCAB06 n009COAXCAB06 n010COAXCAB06 n007COAXCAB06 n008COAXCAB06 1 
R7COAXCAB06 n010COAXCAB06 RBssCOAXCAB06 {Rccoax_2livech} 
E2COAXCAB06 n008COAXCAB06 LBssCOAXCAB06 n010COAXCAB06 RBssCOAXCAB06 1 
R8COAXCAB06 RBssCOAXCAB06 N014 1e-3 
R9COAXCAB06 LBssCOAXCAB06 N007 1e-3 
* <component=coax_2sh>Rs=Rccoax_2shh Ls=Lccoax_2shh RsG=Rccoax_2shg LsG=Lccoax_2shg Cp=Cccoax_2shsh Rp=Rccoax_2shsh k=kccoax_2sh Rch=Rccoax_2shch </component>
.param Rs2_COAXCAB07={0.5*Rccoax_2shh} Ls2_COAXCAB07={0.5*Lccoax_2shh} RsG2_COAXCAB07={0.5*Rccoax_2shg} LsG2_COAXCAB07={0.5*Lccoax_2shg} 
R1COAXCAB07 N031 n001COAXCAB07 {Rs2_COAXCAB07} 
L1COAXCAB07 n001COAXCAB07 n002COAXCAB07 {Ls2_COAXCAB07} 
L2COAXCAB07 n002COAXCAB07 n003COAXCAB07 {Ls2_COAXCAB07} 
R2COAXCAB07 n003COAXCAB07 n007COAXCAB07 {Rs2_COAXCAB07} 
K1COAXCAB07 L1COAXCAB07 L3COAXCAB07 {kccoax_2sh} 
R3COAXCAB07 N013 n004COAXCAB07 {RsG2_COAXCAB07} 
L3COAXCAB07 n004COAXCAB07 n005COAXCAB07 {LsG2_COAXCAB07} 
L4COAXCAB07 n005COAXCAB07 n006COAXCAB07 {LsG2_COAXCAB07} 
R4COAXCAB07 n006COAXCAB07 n009COAXCAB07 {RsG2_COAXCAB07} 
K2COAXCAB07 L2COAXCAB07 L4COAXCAB07 {kccoax_2sh} 
C1COAXCAB07 n002COAXCAB07 n005COAXCAB07 {Cccoax_2shsh} 
R5COAXCAB07 n002COAXCAB07 n005COAXCAB07 {Rccoax_2shsh} 
R6COAXCAB07 n007COAXCAB07 n008COAXCAB07 {Rccoax_2shch} 
E1COAXCAB07 n009COAXCAB07 n010COAXCAB07 n007COAXCAB07 n008COAXCAB07 1 
R7COAXCAB07 n010COAXCAB07 RBssCOAXCAB07 {Rccoax_2shch} 
E2COAXCAB07 n008COAXCAB07 LBssCOAXCAB07 n010COAXCAB07 RBssCOAXCAB07 1 
R8COAXCAB07 RBssCOAXCAB07 N032 1e-3 
R9COAXCAB07 LBssCOAXCAB07 N040 1e-3 
* <twax>\n  Rs={Rs%} Ls={Ls%} RsG={RsG%} LsG={LsG%} Mlg={Mlg%} Cp={Cp%} Rp={Rp%}\n  RsS={RsS%} LsS={LsS%} Mls={Mls%} Mgs={Mgs%} CpS={CpS%} RpS={RpS%}\n  Mll={Mll%} Mgg={Mgg%} Mlg2={Mlg2%} CpGG={CpGG%} RpGG={RpGG%}\n</twax>
* <epbuf>\n  CgA={CgA_%} RgA={RgA_%} CgB={CgB_%} RgB={RgB_%}\n  LoA={LoA_%} RoA={RoA_%} LoB={LoB_%} RoB={RoB_%}\n</epbuf>
* <coax>\n  Rs={Rc%h} Ls={Lc%h} RsG={Rc%g} LsG={Lc%g} Cp={Cc%sh} Rp={Rc%sh} k={kc%} Rch={Rc%ch}\n</coax>
* <adc>\n  Ci={Ca%in} Ri={Ra%in} Clg={Ca%lg} Rlg={Ra%lg} Cgs={Ca%gs} Rgs={Ra%gs} guard={grda%}\n</adc>
* <lug>\n  Ls={R%} Rs={L%}\n</lug>


*** CONTENT OF LIB FILE: E:\smaslan\LV_prog\open-z-bridge-master\sim\ZbrgLib.cir ***
* Twinax cable (two separately shielded cores and one shiled around both)
.SUBCKT TWAXSH AL1 AG1 BL1 BG1 SH1 AL2 AG2 BL2 BG2 SH2 Rs=0.07 Ls=1.1e-6 RsG=0.03 LsG=800e-9 Mlg=790e-9 Cp=95e-12 Rp=1e9 RsS=0.007 LsS=560e-9 Mls=560e-9 Mgs=560e-9 CpS=37e-12 RpS=1e9 Mll=190e-9 Mgg=530e-9 Mlg2=530e-9 CpGG=60e-12 RpGG=1e9
.param Rs2={0.5*Rs} Ls2={0.5*Ls} RsG2={0.5*RsG} LsG2={0.5*LsG} RsS2={0.5*RsS} LsS2={0.5*LsS}
.param Rnull=1e9 $ safety shunts at ends of cables to prevent div by zero when not connected
.param k_lg={Mlg/sqrt(Ls*LsG)} k_ls={Mls/sqrt(Ls*LsS)} k_gs={Mgs/sqrt(LsG*LsS)} k_gg={Mgg/sqrt(LsG*LsG)} k_ll={Mll/sqrt(Ls*Ls)} k_lg2={Mlg2/sqrt(Ls*LsG)}
L1 N003 P001 {LsG2} $ <Lbr> - Cable B return (stray coupling injection point)
L2 N004 P002 {Ls2} $ <Lb> - Cable B live (stray coupling injection point)
L3 P003 N003 {LsG2} $ <Lbr2> - Cable B return (stray coupling injection point)
L4 P004 N004 {Ls2} $ <Lb2> - Cable B live (stray coupling injection point)
C1 N003 N004 {Cp}
R1 N003 N004 {Rp}
R2 P001 BG1 {RsG2}
R3 P002 BL1 {Rs2}
R4 BL2 P004 {Rs2}
R5 BG2 P003 {RsG2}
L5 N001 P005 {Ls2} $ <La> - Cable A live (stray coupling injection point)
L6 N002 P006 {LsG2} $ <Lar> - Cable A return (stray coupling injection point)
L7 P007 N001 {Ls2} $ <La2> - Cable A live (stray coupling injection point)
L8 P008 N002 {LsG2} $ <Lar2> - Cable A return (stray coupling injection point)
C2 N001 N002 {Cp}
R6 N001 N002 {Rp}
R7 P005 AL1 {Rs2}
R8 P006 AG1 {RsG2}
R9 AG2 P008 {RsG2}
R10 AL2 P007 {Rs2}
L9 CAP P009 {LsS2} $ <Lsh> - Outer shield (stray coupling injection point)
L10 P010 CAP {LsS2} $ <Lsh2> - Outer shield (stray coupling injection point)
R11 P009 SH1 {RsS2}
R12 SH2 P010 {RsS2}
C3 N002 CAP {CpS} $ <C:2> - Stray capacitive coupling injection point (format <C:node_id_one_based>)
C4 CAP N003 {CpS}
R13 CAP N003 {RpS}
R14 N002 CAP {RpS}
C5 N002 N003 {CpGG}
R15 N002 N003 {RpGG}
R16 AL1 AG1 {Rnull}
R17 AG1 SH1 {Rnull}
R18 SH1 BG1 {Rnull}
R19 BG1 BL1 {Rnull}
R20 BG2 BL2 {Rnull}
R21 SH2 BG2 {Rnull}
R22 AG2 SH2 {Rnull}
R23 AL2 AG2 {Rnull}
Kla L5 L6 {k_lg}
Kra L7 L8 {k_lg}
Klb L1 L2 {k_lg}
Krb L3 L4 {k_lg}
Kllsa L5 L9 {k_ls}
Klgsa L6 L9 {k_gs}
Klgsb L1 L9 {k_gs}
Kllsb L2 L9 {k_ls}
Klgg L6 L1 {k_gg}
Klll L5 L2 {k_ll}
Klgl L6 L2 {k_lg2}
Klgl2 L5 L1 {k_lg2}
Krlsa L7 L10 {k_ls}
Krgsa L8 L10 {k_gs}
Krgsb L3 L10 {k_gs}
Krlsb L4 L10 {k_ls}
Krgg L8 L3 {k_gg}
Krll L7 L4 {k_ll}
Krgl L8 L4 {k_lg2}
Krgl2 L7 L3 {k_lg2}
.ENDS TWAXSH

* Pair of guard buffers for coax-shields of two cables (twinax cable guard)
.SUBCKT DUAL_EPBUF AL1 AG1 BL1 BG1 AL2 AG2 BL2 BG2 CASE CgA=1e-15 RgA=1e9 CgB=1e-15 RgB=1e9 LoA=1e-12 RoA=1e-6 LoB=1e-12 RoB=1e-6
* cable A
R1 AL1 ep_in_A 1e-3
R2 AL2 ep_in_A 1e-3
R3 AG1 ep_out_A 1e-3
R4 AG2 ep_out_A 1e-3
* buffer A
R11 ep_in_A CASE {RgA}
C1 ep_in_A CASE {CgA}
E1 ep_A1 CASE ep_in_A CASE 1
R5 ep_A1 ep_A2 {RoA}
L1 ep_A2 ep_out_A {LoA}
* cable B
R6 BL1 ep_in_B 1e-3
R7 BL2 ep_in_B 1e-3
R8 BG1 ep_out_B 1e-3
R9 BG2 ep_out_B 1e-3
* buffer B
R12 ep_in_B CASE {RgB}
C2 ep_in_B CASE {CgB}
E2 ep_B1 CASE ep_in_B CASE 1
R10 ep_B1 ep_B2 {RoB}
L2 ep_B2 ep_out_B {LoB}
.ENDS DUAL_EPBUF

* digitizer 3458A with buffered 'isolated' output and internal strays
* optional guarding when 'guard=0' means Rgs||Cgs is ignored and external pin GRD is not connected
.SUBCKT DIG3458 HI LO GRD CASE OUTP OUTN Ci=270e-12 Ri=1e9 Clg=1e-9 Rlg=1e9 Cgs=1e-9 Rgs=1e9 guard=0
* external GRD pin connection only in guarding mode
Rgrd GRD GRDint {(guard>0.5)?1e-6:1e9}
R1 HI LO {Ri}
C1 HI LO {Ci}
E1 OUTP OUTN HI LO 1
R4 LO GRDint {Rlg}
C2 LO GRDint {Clg}
* internal GRD to CASE bridge only in non-guarding mode
R5 GRDint CASE {(guard<0.5)?1e-6:Rgs}
C3 GRDint CASE {Cgs}
R6 OUTP OUTN 1e6
R7 OUTN CASE 1e9
.ENDS DIG3458

* Coax cable with choke having real component
.SUBCKT COAXCAB LA LB RA RB Rs=0.05 Ls=250e-9 RsG=0.05 LsG=250e-9 k=0.9 Cp=105e-12 Rp=1e9 Rch=1e-9
.param Rs2={0.5*Rs} Ls2={0.5*Ls} RsG2={0.5*RsG} LsG2={0.5*LsG}
* high wire
R1 LA n001 {Rs2}
L1 n001 n002 {Ls2} $ <L> - high side tag for inductor for parasitic coupling simulation
L2 n002 n003 {Ls2} $ <L2> - high side tag for inductor for parasitic coupling simulation
R2 n003 n007 {Rs2}
K1 L1 L3 {k}
* low wire
R3 RA n004 {RsG2}
L3 n004 n005 {LsG2} $ <Lg> - low side tag for inductor for parasitic coupling simulation
L4 n005 n006 {LsG2} $ <Lg2> - low side tag for inductor for parasitic coupling simulation
R4 n006 n009 {RsG2}
K2 L2 L4 {k}
* shunting Y
C1 n002 n005 {Cp} $ <C:2> - node tag for capacitor for parasitic coupling simulation
R5 n002 n005 {Rp}
* choke real component simulated
R6 n007 n008 {Rch}
E1 n009 n010 n007 n008 1
R7 n010 RBss {Rch}
E2 n008 LBss n010 RBss 1
R8 RBss RB 1e-3 $ <sense>
R9 LBss LB 1e-3 $ <sense>
* R10 n007 LB 1e-6
* R11 n009 RB 1e-6
.ENDS COAXCAB

* Coax cable with choke having real component and wrapped around wire
.SUBCKT COAXCABGL LA LB RA RB GA GB Rs=0.05 Ls=250e-9 RsR=0.05 LsR=250e-9 k=0.9 Cp=105e-12 Rp=1e9 Rch=1e-9 RsG=0.01 LsG=250e-9 CpG=105e-12 kG=0.9
.param Rs2={0.5*Rs} Ls2={0.5*Ls} RsR2={0.5*RsR} LsR2={0.5*LsR} RsG2={0.5*RsG} LsG2={0.5*LsG}
* high wire
R1 LA n001 {Rs2}
L1 n001 n002 {Ls2} $ <L> - high side tag for inductor for parasitic coupling simulation
L2 n002 n003 {Ls2} $ <L2> - high side tag for inductor for parasitic coupling simulation
R2 n003 n007 {Rs2}
K1 L1 L3 {k}
* low wire
R3 RA n004 {RsR2}
L3 n004 n005 {LsR2} $ <Lr> - low side tag for inductor for parasitic coupling simulation
L4 n005 n006 {LsR2} $ <Lr2> - low side tag for inductor for parasitic coupling simulation
R4 n006 n009 {RsR2}
K2 L2 L4 {k}
* shunting Y
C1 n002 n005 {Cp} $ <C:2> - node tag for capacitor for parasitic coupling simulation
R5 n002 n005 {Rp}
* choke real component simulated
R6 n007 n008 {Rch}
E1 n009 n010 n007 n008 1
R7 n010 RBss {Rch}
E2 n008 LBss n010 RBss 1
* auxiliary wire
Rw1 GA w001 {RsG2}
Lw1 w001 w002 {LsG2} $ <Lg> - gnd lug coupling
Lw2 w002 w003 {LsG2} $ <Lg2> - gnd lug coupling
Rw2 w003 GBss {RsG2}
Cw w002 n005 {CpG} $ <C:1> - capacitive coupling to ground lug
K3 L1 Lw1 {kG}
K4 L3 Lw1 {kG}
K5 L2 Lw2 {kG}
K6 L4 Lw2 {kG}
* current sensing
R8 RBss RB 1e-3 $ <sense>
R9 LBss LB 1e-3 $ <sense>
R10 GBss GB 1e-3 $ <sense>
.ENDS COAXCABGL

* Coax cable
.SUBCKT COAXCAB2 LA LB RA RB Rs=0.05 Ls=250e-9 RsG=0.05 LsG=250e-9 k=0.9 Cp=105e-12 Rp=1e9
R1 LA n001 {Rs}
L1 n001 n002 {Ls}
L2 n002 n003 {Ls}
R2 n003 LB {Rs}
R3 RA n004 {RsG}
L3 n004 n005 {LsG}
L4 n005 n006 {LsG}
R4 n006 RB {RsG}
C1 n002 n005 {Cp}
R5 n002 n005 {Rp}
K1 L1 L3 {k}
K2 L2 L4 {k}
.ENDS COAXCAB2

* Ground lug
.SUBCKT GNDLUG LA LB Rs=0.05 Ls=250e-9
R1 LA n001 {Rs} $ <C:2> - capacitance injection point
L1 n001 LB {Ls} $ <L> - high side tag for inductor for parasitic coupling simulation
.ENDS GNDLUG

* 4TP standard
.SUBCKT STD4TP Hp HpG Lp LpG Hc HcG Lc LcG COM Rp=0.01 Lp=20e-9 Rpg=0.005 Lpg=15e-9 kp=0.7 Cps=5e-12 Rps=1e9 Rc=0.01 Lc=20e-9 Rcg=0.005 Lcg=15e-9 kc=0.7 Ccs=5e-12 Rcs=1e9 Rs=100 Ls=0
R1 high n001 {Rs}
L1 n001 low {Ls}
Xhpot Hp high HpG COM COAXCAB2 Rs={Rp} Ls={Lp} RsG={Rpg} LsG={Lpg} k={kp} Cp={Cps} Rp={Rps}
Xlpot Lp low LpG COM COAXCAB2 Rs={Rp} Ls={Lp} RsG={Rpg} LsG={Lpg} k={kp} Cp={Cps} Rp={Rps}
Xhcur Hc high HcG COM COAXCAB2 Rs={Rc} Ls={Lc} RsG={Rcg} LsG={Lcg} k={kc} Cp={Ccs} Rp={Rcs}
Xlcur Lc low LcG COM COAXCAB2 Rs={Rc} Ls={Lc} RsG={Rcg} LsG={Lcg} k={kc} Cp={Ccs} Rp={Rcs}
.ENDS STD4TP

* 4TP standard with split grounds
.SUBCKT STD4TP2 Hp HpG Lp LpG Hc HcG Lc LcG Gp Gc Rp=0.01 Lp=20e-9 Rpg=0.005 Lpg=15e-9 kp=0.7 Cps=5e-12 Rps=1e9 Rc=0.01 Lc=20e-9 Rcg=0.005 Lcg=15e-9 kc=0.7 Ccs=5e-12 Rcs=1e9 Rs=100 Ls=0
R1 high n001 {Rs}
L1 n001 low {Ls}
Xhpot Hp high HpG Gp COAXCAB2 Rs={Rp} Ls={Lp} RsG={Rpg} LsG={Lpg} k={kp} Cp={Cps} Rp={Rps}
Xlpot Lp low LpG Gp COAXCAB2 Rs={Rp} Ls={Lp} RsG={Rpg} LsG={Lpg} k={kp} Cp={Cps} Rp={Rps}
Xhcur Hc high HcG Gc COAXCAB2 Rs={Rc} Ls={Lc} RsG={Rcg} LsG={Lcg} k={kc} Cp={Ccs} Rp={Rcs}
Xlcur Lc low LcG Gc COAXCAB2 Rs={Rc} Ls={Lc} RsG={Rcg} LsG={Lcg} k={kc} Cp={Ccs} Rp={Rcs}
.ENDS STD4TP2

* realistic 4TP standard with optional split grounds and optional return path impedance
.SUBCKT STD4TP3 Hp HpG Lp LpG Hc HcG Lc LcG Gp Gc Rp=0.01 Lp=20e-9 Rpg=0.005 Lpg=15e-9 kp=0.7 Cps=5e-12 Rps=1e9 Rc=0.01 Lc=20e-9 Rcg=0.005 Lcg=15e-9 kc=0.7 Ccs=5e-12 Rcs=1e9 Rs=100 Ls=0 Rg=1e-11 Lg=1 Rb=1e-11 Lb=1
.param Rgx={(abs(Rg)>5e-10)?Rg:1e-9} Lgx={(abs(Rg)>5e-10)?Lg:1e-12} Rpg1={(abs(Rg)>5e-10)?1e9:1e-9} Rpg2={(abs(Rg)>5e-10)?1e-9:1e9}
.param Rcg1={(abs(Rg)>5e-10)?1e9:1e-9} Rcg2=1e-9 Rcg3={(abs(Rg)>5e-10)?1e9:1e-9}
L1 N006 N010 {Ls}
R1 N001 N006 {Rs}
R2 N003 N002 {Rb}
L2 N004 N003 {Lb}
R3 N009 N008 {Rb}
L3 N007 N009 {Lb}
R4 P001 N002 {0.5*Rgx}
L4 N005 P001 {0.5*Lgx}
R5 P002 N008 {0.5*Rgx}
L5 N005 P002 {0.5*Lgx}
R6 N007 N004 {Rcg1}
R7 N004 Gc {Rcg2}
R8 N007 Gc {Rcg3}
R9 Gp N005 {Rpg1}
R10 Gp N002 {Rpg2}
XHC Hc N001 HcG N004 COAXCAB2 Rs={Rc} Ls={Lc} RsG={Rcg} LsG={Lcg} k={kc} Cp={Ccs} Rp={Rcs}
XLC N010 Lc N007 LcG COAXCAB2 Rs={Rc} Ls={Lc} RsG={Rcg} LsG={Lcg} k={kc} Cp={Ccs} Rp={Rcs}
XHP Hp N001 HpG N002 COAXCAB2 Rs={Rp} Ls={Lp} RsG={Rpg} LsG={Lpg} k={kp} Cp={Cps} Rp={Rps}
XLP Lp N010 LpG N008 COAXCAB2 Rs={Rp} Ls={Lp} RsG={Rpg} LsG={Lpg} k={kp} Cp={Cps} Rp={Rps}
.ENDS STD4TP3

* Coaxial standard
.SUBCKT STDCOAX Ch Cl Ph Pl Rp=0.01 Lp=20e-9 Rpg=0.005 Lpg=15e-9 kp=0.7 Cps=5e-12 Rps=1e9 Rc=0.01 Lc=20e-9 Rcg=0.005 Lcg=15e-9 kc=0.7 Ccs=5e-12 Rcs=1e9 Rs=1 Ls=0
R1 high n001 {Rs}
L1 n001 low {Ls}
Xcur Ch high Cl low COAXCAB2 Rs={Rc} Ls={Lc} RsG={Rcg} LsG={Lcg} k={kc} Cp={Ccs} Rp={Rcs}
Xpot Ph high Pl low COAXCAB2 Rs={Rp} Ls={Lp} RsG={Rpg} LsG={Lpg} k={kp} Cp={Cps} Rp={Rps}
.ENDS STDCOAX

* Coaxial standard with 2x2TP adapters (4TP)
.SUBCKT STDCOAX4TP Ch ChG Cl ClG Ph PhG Pl PlG Rp=0.01 Lp=20e-9 Rpg=0.005 Lpg=15e-9 kp=0.7 Cps=5e-12 Rps=1e9 Rc=0.01 Lc=20e-9 Rcg=0.005 Lcg=15e-9 kc=0.7 Ccs=5e-12 Rcs=1e9 Rs=1 Ls=0
* shunt impedance
R1 high n001 {Rs}
L1 n001 low {Ls}
* current ports
XcurH Ch high ChG Cgnd1 COAXCAB2 Rs={Rc} Ls={Lc} RsG={Rcg} LsG={Lcg} k={kc} Cp={Ccs} Rp={Rcs}
XcurL Cl low ClG Cgnd2 COAXCAB2 Rs={Rc} Ls={Lc} RsG={Rcg} LsG={Lcg} k={kc} Cp={Ccs} Rp={Rcs}
R2 Cgnd1 Cgnd2 0.0001
* potential ports
XpotH Ph high PhG Pgnd1 COAXCAB2 Rs={Rp} Ls={Lp} RsG={Rpg} LsG={Lpg} k={kp} Cp={Cps} Rp={Rps}
XpotL Pl low PlG Pgnd2 COAXCAB2 Rs={Rp} Ls={Lp} RsG={Rpg} LsG={Lpg} k={kp} Cp={Cps} Rp={Rps}
R3 Pgnd1 Pgnd2 0.0001
.ENDS STDCOAX4TP

* Coaxial standard with 1P input and 2TP output
.SUBCKT STDCOAX1P2TP Ch Cl Ph PhG Pl PlG Rp=0.01 Lp=20e-9 Rpg=0.005 Lpg=15e-9 kp=0.7 Cps=5e-12 Rps=1e9 Rc=0.01 Lc=20e-9 Rcg=0.005 Lcg=15e-9 kc=0.7 Ccs=5e-12 Rcs=1e9 Rs=1 Ls=0
* shunt impedance
R1 high n001 {Rs}
L1 n001 low {Ls}
* current ports
XcurH Ch high Cl low COAXCAB2 Rs={Rc} Ls={Lc} RsG={Rcg} LsG={Lcg} k={kc} Cp={Ccs} Rp={Rcs}
* potential ports
XpotH Ph high PhG Pgnd1 COAXCAB2 Rs={Rp} Ls={Lp} RsG={Rpg} LsG={Lpg} k={kp} Cp={Cps} Rp={Rps}
XpotL Pl low PlG Pgnd2 COAXCAB2 Rs={Rp} Ls={Lp} RsG={Rpg} LsG={Lpg} k={kp} Cp={Cps} Rp={Rps}
R2 Pgnd1 Pgnd2 0.0001
.ENDS STDCOAX1P2TP



* LF 4TP Kelvin injection transformer
* Lp-Rp-Cp: primary
* Ls-Rs: secondary
* k: coupling
* ksh: shields half-turn coupling
* Lsh-Rsh: shield half-loop impedance
* Csl1, Csl2: shield 1 and 2 loop capacitance
* C12a,b: primary to shield 1 capacitances (Z1-a, Z2-b)
* C23a,b: shield 1 to shield 2 capacitances (Z1-a, Z2-b)
* C34a,b: shield 2 to shield secondary capacitances (Z1-a, Z2-b)
.SUBCKT LF4TPKETR Z1 Z1G Z2 Z2G IN1 IN2 SH1 SH2 Lp=1 Rp=1 Cp=100e-12 Ls=10e-6 Rs=0.001 k=0.999 ksh=0.999 Lsh=2.5e-6 Rsh=1 Csl1=5e-12 Csl2=5e-12 C12a=100e-12 C12b=100e-12 C23a=100e-12 C23b=100e-12 C34a=100e-12 C34b=100e-12
L1 IN1 P001 {Lp}
L2 Z1 P002 {Ls}
L3 N001 N003 {Lsh}
L4 N005 N007 {Lsh}
C1 N003 N005 {Csl1}
C2 IN1 IN2 {Cp}
C3 N003 P003 {C12a}
C4 N005 P004 {C12b}
L5 N002 N004 {Lsh}
L6 N006 N008 {Lsh}
C5 N004 N006 {Csl2}
C6 N004 P005 {C23a}
C7 N006 P006 {C23b}
C8 Z1 P007 {C34a}
C9 Z2 P008 {C34b}
R1 P002 Z2 {Rs}
R2 P001 IN2 {Rp}
R3 N001 SH1 {Rsh}
R4 N007 SH1 {Rsh}
R5 Z2G N008 {Rsh}
R6 Z1G N002 {Rsh}
R7 P005 N003 1
R8 P006 N005 1
R9 P003 IN1 1
R10 P004 IN2 1
R11 P007 N004 1
R12 P008 N006 1
R13 Z1G SH2 1e-3
R14 SH2 Z2G 1e-3
K1 L1 L2 {k}
K2 L1 L3 {ksh}
K3 L1 L4 {ksh}
K6 L1 L5 {ksh}
K7 L1 L6 {ksh}
K4 L2 L3 {ksh}
K5 L2 L4 {ksh}
K8 L2 L5 {ksh}
K9 L2 L6 {ksh}
.ENDS LF4TPKETR


* LF coaxial Kelvin injection transformer
* Lp-Rp-Cp: primary
* Ls-Rs: secondary
* k: coupling
* ksh: shields half-turn coupling
* Lsh-Rsh: shield half-loop impedance
* Csl1, Csl2: shield 1 and 2 loop capacitance
* C12a,b: primary to shield 1 capacitances (Z1-a, Z2-b)
* C23a,b: shield 1 to shield 2 capacitances (Z1-a, Z2-b)
* C34a,b: shield 2 to shield secondary capacitances (Z1-a, Z2-b)
* C45a,b: secondary to main supply capacitances (Z1-a, Z2-b)
.SUBCKT LFCOAXKETR Z1 Z1G Z2 Z2G IN1 IN2 M1 M2 SH1 SH2 Lp=1 Rp=1 Cp=100e-12 Ls=10e-6 Rs=0.001 k=0.999 ksh=0.999 Lsh=2.5e-6 Rsh=1 Csl1=5e-12 Csl2=5e-12 C12a=100e-12 C12b=100e-12 C23a=100e-12 C23b=100e-12 C34a=100e-12 C34b=100e-12 C45a=100e-12 C45b=100e-12
L1 IN1 P001 {Lp}
L2 Z1G P002 {Ls}
L3 N001 N003 {Lsh}
L4 N005 N007 {Lsh}
C1 N003 N005 {Csl1}
C2 IN1 IN2 {Cp}
C3 N003 P003 {C12a}
C4 N005 P004 {C12b}
L5 N002 N004 {Lsh}
L6 N006 N008 {Lsh}
C5 N004 N006 {Csl2}
C6 N004 P005 {C23a}
C7 N006 P006 {C23b}
C8 Z1G P007 {C34a}
C9 Z2G P008 {C34b}
R1 P002 Z2G {Rs}
C10 M1 SH2 {C45a}
C11 M2 SH2 {C45b}
R2 P001 IN2 {Rp}
R3 N001 SH1 {Rsh}
R4 N007 SH1 {Rsh}
R5 SH2 N008 {Rsh}
R6 SH2 N002 {Rsh}
R7 P005 N003 1
R8 P006 N005 1
R9 P003 IN1 1
R10 P004 IN2 1
R11 P007 N004 1
R12 P008 N006 1
R13 Z1 M1 1e-6
R14 M2 Z2 1e-6
K1 L1 L2 {k}
K2 L1 L3 {ksh}
K3 L1 L4 {ksh}
K6 L1 L5 {ksh}
K7 L1 L6 {ksh}
K4 L2 L3 {ksh}
K5 L2 L4 {ksh}
K8 L2 L5 {ksh}
K9 L2 L6 {ksh}
.ENDS LFCOAXKETR

* LF main transformer
*  Lp-Rp-Cp: primary
*  Ls-Rs: secondary
*  k: coupling
*  ksh: shields half-turn coupling
*  Lsh-Rsh: shield half-loop impedance
*  Csl1, Csl2: shield 1 and 2 loop capacitance
*  C12a,b: primary to shield 1 capacitances (Z1-a, Z2-b)
*  C23a,b: shield 1 to shield 2 capacitances (Z1-a, Z2-b)
*  C34a,b: shield 2 to shield secondary capacitances (Z1-a, Z2-b)
.SUBCKT LFMAINTR IN1 IN2 SH1 OUT1 OUT2 SH2 Lp=1 Rp=1 Cp=100e-12 Ls=10e-6 Rs=0.001 k=0.999 ksh=0.999 Lsh=2.5e-6 Rsh=1 Csl1=5e-12 Csl2=5e-12 C12a=100e-12 C12b=100e-12 C23a=100e-12 C23b=100e-12 C34a=100e-12 C34b=100e-12
L1 IN1 P001 {Lp}
L2 OUT1 P002 {Ls}
L3 N001 UR1 {Lsh}
L4 UR2 N005 {Lsh}
C1 UR1 UR2 {Csl1}
C2 IN1 IN2 {Cp}
C3 UR1 P003 {C12a}
C4 UR2 P004 {C12b}
L5 N002 N003 {Lsh}
L6 N004 N006 {Lsh}
C5 N003 N004 {Csl2}
C6 N003 P005 {C23a}
C7 N004 P006 {C23b}
C8 OUT1 P007 {C34a}
C9 OUT2 P008 {C34b}
R1 P002 OUT2 {Rs}
R2 P001 IN2 {Rp}
R3 N001 SH1 {Rsh}
R4 N005 SH1 {Rsh}
R5 SH2 N006 {Rsh}
R6 SH2 N002 {Rsh}
R7 P005 UR1 1
R8 P006 UR2 1
R9 P003 IN1 1
R10 P004 IN2 1
R11 P007 N003 1
R12 P008 N004 1
K1 L1 L2 {k}
K2 L1 L3 {ksh}
K3 L1 L4 {ksh}
K6 L1 L5 {ksh}
K7 L1 L6 {ksh}
K4 L2 L3 {ksh}
K5 L2 L4 {ksh}
K8 L2 L5 {ksh}
K9 L2 L6 {ksh}
.ENDS LFMAINTR

* LF main transformer with 3 shields
*  Lp-Rp-Cp: primary
*  Ls-Rs: secondary
*  k: coupling
*  ksh: shields half-turn coupling (must be ksh<k to keep system positive definite)
*  Lsh-Rsh: shield half-loop impedance
*  Csl1, Csl2: shield 1 and 2 loop capacitance
*  C12a,b: primary to shield 1 capacitances (Z1-a, Z2-b)
*  C23a,b: shield 1 to shield 2 capacitances (Z1-a, Z2-b)
*  C34a,b: shield 2 to shield 3 capacitances (Z1-a, Z2-b)
*  C45a,b: shield 3 to shield secondary capacitances (Z1-a, Z2-b)
.SUBCKT LFMAINTR3 IN1 IN2 SH1 OUT1 OUT2 SH2 SH3 Lp=1 Rp=1 Cp=100e-12 Ls=10e-6 Rs=0.001 k=0.999 ksh=0.999 Lsh=2.5e-6 Rsh=1 Csl1=5e-12 Csl2=5e-12 Csl3=5e-12 C12a=100e-12 C12b=100e-12 C23a=100e-12 C23b=100e-12 C34a=100e-12 C34b=100e-12 C45a=100e-12 C45b=100e-12
L1 IN1 P001 {Lp}
L2 OUT1 P002 {Ls}
L3 N001 UR1 {Lsh}
L4 UR2 N008 {Lsh}
C1 UR1 UR2 {Csl1}
C2 IN1 IN2 {Cp}
C3 UR1 P003 {C12a}
C4 UR2 P004 {C12b}
L5 N002 N005 {Lsh}
L6 N007 N010 {Lsh}
C5 N005 N007 {Csl3}
C6 N004 P005 {C23a}
C7 N006 P006 {C23b}
C8 OUT1 P007 {C45a}
C9 OUT2 P008 {C45b}
R1 P002 OUT2 {Rs}
R2 P001 IN2 {Rp}
R3 N001 SH1 {Rsh}
R4 N008 SH1 {Rsh}
R5 SH2 N010 {Rsh}
R6 SH2 N002 {Rsh}
R7 P005 UR1 1
R8 P006 UR2 1
R9 P003 IN1 1
R10 P004 IN2 1
R11 P007 N005 1
R12 P008 N007 1
L7 N003 N004 {Lsh}
L8 N006 N009 {Lsh}
C10 N005 P009 {C34a}
C11 N007 P010 {C34b}
R13 P009 N004 1
R14 P010 N006 1
C12 N004 N006 {Csl2}
R15 N003 SH3 {Rsh}
R16 SH3 N009 {Rsh}
K1 L1 L2 {k}
K2 L1 L3 {ksh}
K3 L1 L4 {ksh}
K9 L2 L3 {ksh}
K10 L2 L4 {ksh}
K4 L1 L5 {ksh}
K5 L1 L6 {ksh}
K11 L2 L5 {ksh}
K12 L2 L6 {ksh}
K7 L1 L7 {ksh}
K8 L1 L8 {ksh}
K13 L2 L7 {ksh}
K14 L2 L8 {ksh}
.ENDS LFMAINTR3

* Twisted cable with shield
.SUBCKT TWCABSH A1 B1 SH1 A2 B2 SH2 Rsa=0.001 Lsa=100e-9 Rsb=0.001 Lsb=100e-9 Cab=50e-12 Cag=20e-12 Cbg=20e-12 k=0.9
.param Rsa2={0.5*Rsa} Rsb2={0.5*Rsb} Lsa2={0.5*Lsa} Lsb2={0.5*Lsb}
R1 N001 A1 {Rsa2}
R2 A2 N003 {Rsa2}
R3 N005 B1 {Rsb2}
R4 B2 N007 {Rsb2}
L1 N001 N002 {Lsa2} $ <L1>
L2 N002 N003 {Lsa2} $ <L2>
L3 N005 N006 {Lsb2} $ <L3>
L4 N006 N007 {Lsb2} $ <L4>
C1 N002 N006 {Cab}
C2 N002 N004 {Cag}
C3 N004 N006 {Cbg}
R5 N004 SH1 1e-3
R6 SH2 N004 1e-3
K1 L1 L3 {k}
K2 L2 L4 {k}
.ENDS TWCABSH

* common mode detector for coaxial cable:
*  Ld: detector inductance
*  n: detector turns count
*  k: coupling
*  Cws: primary winding-shield capacitance (total from both winding ends)
*  Csc: shield-coax capacitance (total to both ends of coax)
.SUBCKT COMDET LA RA LB RB DA DB SH Ld=0.2 n=100 k=0.998 Cws=50e-12 Csc=5e-12
.param Ls={Ld/n^2}
L1 LA LB {Ls}
L2 RA RB {Ls}
L3 DA DB {Ld}
K1 L1 L3 {k}
K2 L2 L3 {k}
K3 L1 L2 {k}
* stray capacitances
Rsh SH SHi 1e-4 $ isolation needed to prevent singular matrix errors
Cws1 DA SHi {0.5*Cws}
Cws2 DB SHi {0.5*Cws}
Csc1 RA SHi {0.5*Csc}
Csc2 RB SHi {0.5*Csc}
.ENDS COMDET

* common mode detector for two coaxial cables:
*  Ld: detector inductance
*  n: detector turns count
*  k: coupling
*  m: mode (0-disabled,1-only to coax 1,2-to both coaxes)
*  Cws: primary winding-shield capacitance (total from both winding ends)
*  Csc1: shield-coax 1 capacitance (total to both ends of coax)
*  Csc2: shield-coax 2 capacitance (total to both ends of coax)
.SUBCKT COMDET2 L1A R1A L1B R1B L2A R2A L2B R2B DA DB SH Ld=0.2 n=100 k=0.998 m=2 Cws=50e-12 Csc1=5e-12 Csc2=5e-12
.param Ls={Ld/n^2}
L1 L1A L1B {(m>0.01)?Ls:1e-9}
L2 R1A R1B {(m>0.01)?Ls:1e-9}
L3 L2A L2B {(m>1.99)?Ls:1e-9}
L4 R2A R2B {(m>1.99)?Ls:1e-9}
L5 DA DB {Ld}
*
K1 L1 L2 {(m>0.01)?k:0.99999}
K2 L1 L3 {(m>1.99)?k:0}
K3 L1 L4 {(m>1.99)?k:0}
K4 L2 L3 {(m>1.99)?k:0}
K5 L2 L4 {(m>1.99)?k:0}
K6 L3 L4 {(m>1.99)?k:0.99999}
*
K7 L5 L1 {(m>0)?k:0}
K8 L5 L2 {(m>0)?k:0}
K9 L5 L3 {(m>1.99)?k:0}
K10 L5 L4 {(m>1.99)?k:0}
* strays
Rsh SH SHi 1e-4 $ isolation needed to prevent singular matrix errors
Cws1 DA SHi {0.5*Cws}
Cws2 DB SHi {0.5*Cws}
Csc1a R1A SHi {(m>0.01)?(0.5*Csc1):1e-15}
Csc1b R1B SHi {(m>0.01)?(0.5*Csc1):1e-15}
Csc2a R2A SHi {(m>1.99)?(0.5*Csc2):1e-15}
Csc2b R2B SHi {(m>1.99)?(0.5*Csc2):1e-15}
.ENDS COMDET2


* buffer with phase shifting
*  g: gain
*  ph: phase shift in [rad] in range (-pi/2:+pi/2) only!
*  Cp-Rp: input shunting
*  Ls-Rs: output impedance
.SUBCKT BUFPHI IN OUT REF g=1 ph=0 Cp=5e-12 Rp=1e6 Rs=0.001 Ls=100e-9
* input shunting
Rin IN REF {Rp}
Cin IN REF {Cp}
* phase shift +-90deg
B90 V90 REF I=v(IN)*hertz*2*pi*((ph<0)?-1:1)
C90 V90 REF 1
R90 V90 REF 1e9
* mix re/im to get desired phase angle
Bout VOUT REF V=(v(IN)*cos(ph)+v(V90)*sin(abs(ph)))*g
* output impedance
Rout VOUT n001 {Rs}
Lout n001 OUT {Ls}
.ENDS BUFPHI

* 4TP standard ground isolator (splits 1 and 2 side grounds, but keeps coaxial connection)
*  Lsa-Rsa: 1-2 side live signal series impedance cable A
*  Lsb-Rsb: 1-2 side live signal series impedance cable B
*  Lg1-Rg1: side 1 A-B coax ground series impedance
*  Lg2-Rg2: side 2 A-B coax ground series impedance
*  Cab: coax A-B live capacitance
*  C12: capacitance between 1-2 side grounds
*  kab: coupling between A-B lives
*  k12: coupling between side 1-2 grounds
*  Rbyp: side 1-2 grounds bypass
.SUBCKT ISOL4TP A2 A2g B2 B2g A1 A1g B1 B1g G1 G2 Lsa=10e-9 Rsa=2e-3 Lsb=10e-9 Rsb=2e-3 Lg1=10e-9 Rg1=0.5e-3 Lg2=15e-9 Rg2=2e-3 Cab=5e-12 C12=1e-15 kab=0.5 k12=0.5 Rbyp=1e9
L1 N001 A2 {0.5*Lsa}
R1 N002 N001 {0.5*Rsa}
L2 N008 B2 {0.5*Lsb}
R2 N009 N008 {0.5*Rsb}
L3 N005 A1g {0.5*Lg1}
R3 G1 N005 {0.5*Rg1}
L4 N004 A2g {0.5*Lg2}
R4 G2 N004 {0.5*Rg2}
L5 N003 A1 {0.5*Lsa}
R5 N002 N003 {0.5*Rsa}
L6 N010 B1 {0.5*Lsb}
R6 N009 N010 {0.5*Rsb}
L7 N007 B1g {0.5*Lg1}
R7 G1 N007 {0.5*Rg1}
L8 N006 B2g {0.5*Lg2}
R8 G2 N006 {0.5*Rg2}
C1 G1 G2 {C12}
C2 N009 N002 {Cab}
R10 A1g A2g {Rbyp}
R9 B1g B2g {Rbyp}
Kab L1 L2 {kab}
K12 L3 L4 {k12}
K12b L7 L8 {k12}
Kab2 L5 L6 {kab}
.ENDS ISOL4TP


*** END OF CONTENT OF LIB FILE: E:\smaslan\LV_prog\open-z-bridge-master\sim\ZbrgLib.cir ***

* Automatically generated stray couplings
Kstray0001 L1TWAXSH01 L1TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)} $ M#001=<M_stray001>
Kstray0002 L1TWAXSH01 L2TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0003 L1TWAXSH01 L3TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0004 L1TWAXSH01 L4TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0005 L1TWAXSH01 L5TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0006 L1TWAXSH01 L6TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0007 L1TWAXSH01 L7TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0008 L1TWAXSH01 L8TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0009 L1TWAXSH01 L9TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0010 L1TWAXSH01 L10TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0011 L2TWAXSH01 L1TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0012 L2TWAXSH01 L2TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0013 L2TWAXSH01 L3TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0014 L2TWAXSH01 L4TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0015 L2TWAXSH01 L5TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0016 L2TWAXSH01 L6TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0017 L2TWAXSH01 L7TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0018 L2TWAXSH01 L8TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0019 L2TWAXSH01 L9TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0020 L2TWAXSH01 L10TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0021 L3TWAXSH01 L1TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0022 L3TWAXSH01 L2TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0023 L3TWAXSH01 L3TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0024 L3TWAXSH01 L4TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0025 L3TWAXSH01 L5TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0026 L3TWAXSH01 L6TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0027 L3TWAXSH01 L7TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0028 L3TWAXSH01 L8TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0029 L3TWAXSH01 L9TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0030 L3TWAXSH01 L10TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0031 L4TWAXSH01 L1TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0032 L4TWAXSH01 L2TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0033 L4TWAXSH01 L3TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0034 L4TWAXSH01 L4TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0035 L4TWAXSH01 L5TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0036 L4TWAXSH01 L6TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0037 L4TWAXSH01 L7TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0038 L4TWAXSH01 L8TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0039 L4TWAXSH01 L9TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0040 L4TWAXSH01 L10TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0041 L5TWAXSH01 L1TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0042 L5TWAXSH01 L2TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0043 L5TWAXSH01 L3TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0044 L5TWAXSH01 L4TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0045 L5TWAXSH01 L5TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0046 L5TWAXSH01 L6TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0047 L5TWAXSH01 L7TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0048 L5TWAXSH01 L8TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0049 L5TWAXSH01 L9TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0050 L5TWAXSH01 L10TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0051 L6TWAXSH01 L1TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0052 L6TWAXSH01 L2TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0053 L6TWAXSH01 L3TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0054 L6TWAXSH01 L4TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0055 L6TWAXSH01 L5TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0056 L6TWAXSH01 L6TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0057 L6TWAXSH01 L7TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0058 L6TWAXSH01 L8TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0059 L6TWAXSH01 L9TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0060 L6TWAXSH01 L10TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0061 L7TWAXSH01 L1TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0062 L7TWAXSH01 L2TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0063 L7TWAXSH01 L3TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0064 L7TWAXSH01 L4TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0065 L7TWAXSH01 L5TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0066 L7TWAXSH01 L6TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0067 L7TWAXSH01 L7TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0068 L7TWAXSH01 L8TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0069 L7TWAXSH01 L9TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0070 L7TWAXSH01 L10TWAXSH02 {max(min(M_stray001/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0071 L8TWAXSH01 L1TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0072 L8TWAXSH01 L2TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0073 L8TWAXSH01 L3TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0074 L8TWAXSH01 L4TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0075 L8TWAXSH01 L5TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0076 L8TWAXSH01 L6TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0077 L8TWAXSH01 L7TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0078 L8TWAXSH01 L8TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0079 L8TWAXSH01 L9TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0080 L8TWAXSH01 L10TWAXSH02 {max(min(M_stray001/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0081 L9TWAXSH01 L1TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0082 L9TWAXSH01 L2TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0083 L9TWAXSH01 L3TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0084 L9TWAXSH01 L4TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0085 L9TWAXSH01 L5TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0086 L9TWAXSH01 L6TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0087 L9TWAXSH01 L7TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0088 L9TWAXSH01 L8TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0089 L9TWAXSH01 L9TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0090 L9TWAXSH01 L10TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0091 L10TWAXSH01 L1TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0092 L10TWAXSH01 L2TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0093 L10TWAXSH01 L3TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0094 L10TWAXSH01 L4TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0095 L10TWAXSH01 L5TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0096 L10TWAXSH01 L6TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0097 L10TWAXSH01 L7TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray0098 L10TWAXSH01 L8TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray0099 L10TWAXSH01 L9TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray0100 L10TWAXSH01 L10TWAXSH02 {max(min(M_stray001/sqrt(abs(LsS2_TWAXSH01*LsS2_TWAXSH02)),0.999),-0.999)}
Cstray001 CAPTWAXSH01 CAPTWAXSH02 {C_stray001} $ C#001=<C_stray001>
Kstray0101 L1TWAXSH03 L1TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)} $ M#002=<M_stray002>
Kstray0102 L1TWAXSH03 L2TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0103 L1TWAXSH03 L3TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0104 L1TWAXSH03 L4TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0105 L1TWAXSH03 L5TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0106 L1TWAXSH03 L6TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0107 L1TWAXSH03 L7TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0108 L1TWAXSH03 L8TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0109 L1TWAXSH03 L9TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0110 L1TWAXSH03 L10TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0111 L2TWAXSH03 L1TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0112 L2TWAXSH03 L2TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0113 L2TWAXSH03 L3TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0114 L2TWAXSH03 L4TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0115 L2TWAXSH03 L5TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0116 L2TWAXSH03 L6TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0117 L2TWAXSH03 L7TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0118 L2TWAXSH03 L8TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0119 L2TWAXSH03 L9TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0120 L2TWAXSH03 L10TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0121 L3TWAXSH03 L1TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0122 L3TWAXSH03 L2TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0123 L3TWAXSH03 L3TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0124 L3TWAXSH03 L4TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0125 L3TWAXSH03 L5TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0126 L3TWAXSH03 L6TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0127 L3TWAXSH03 L7TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0128 L3TWAXSH03 L8TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0129 L3TWAXSH03 L9TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0130 L3TWAXSH03 L10TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0131 L4TWAXSH03 L1TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0132 L4TWAXSH03 L2TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0133 L4TWAXSH03 L3TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0134 L4TWAXSH03 L4TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0135 L4TWAXSH03 L5TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0136 L4TWAXSH03 L6TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0137 L4TWAXSH03 L7TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0138 L4TWAXSH03 L8TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0139 L4TWAXSH03 L9TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0140 L4TWAXSH03 L10TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0141 L5TWAXSH03 L1TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0142 L5TWAXSH03 L2TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0143 L5TWAXSH03 L3TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0144 L5TWAXSH03 L4TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0145 L5TWAXSH03 L5TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0146 L5TWAXSH03 L6TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0147 L5TWAXSH03 L7TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0148 L5TWAXSH03 L8TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0149 L5TWAXSH03 L9TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0150 L5TWAXSH03 L10TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0151 L6TWAXSH03 L1TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0152 L6TWAXSH03 L2TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0153 L6TWAXSH03 L3TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0154 L6TWAXSH03 L4TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0155 L6TWAXSH03 L5TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0156 L6TWAXSH03 L6TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0157 L6TWAXSH03 L7TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0158 L6TWAXSH03 L8TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0159 L6TWAXSH03 L9TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0160 L6TWAXSH03 L10TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0161 L7TWAXSH03 L1TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0162 L7TWAXSH03 L2TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0163 L7TWAXSH03 L3TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0164 L7TWAXSH03 L4TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0165 L7TWAXSH03 L5TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0166 L7TWAXSH03 L6TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0167 L7TWAXSH03 L7TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0168 L7TWAXSH03 L8TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0169 L7TWAXSH03 L9TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0170 L7TWAXSH03 L10TWAXSH04 {max(min(M_stray002/sqrt(abs(Ls2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0171 L8TWAXSH03 L1TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0172 L8TWAXSH03 L2TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0173 L8TWAXSH03 L3TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0174 L8TWAXSH03 L4TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0175 L8TWAXSH03 L5TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0176 L8TWAXSH03 L6TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0177 L8TWAXSH03 L7TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0178 L8TWAXSH03 L8TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0179 L8TWAXSH03 L9TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0180 L8TWAXSH03 L10TWAXSH04 {max(min(M_stray002/sqrt(abs(LsG2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0181 L9TWAXSH03 L1TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0182 L9TWAXSH03 L2TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0183 L9TWAXSH03 L3TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0184 L9TWAXSH03 L4TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0185 L9TWAXSH03 L5TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0186 L9TWAXSH03 L6TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0187 L9TWAXSH03 L7TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0188 L9TWAXSH03 L8TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0189 L9TWAXSH03 L9TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0190 L9TWAXSH03 L10TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0191 L10TWAXSH03 L1TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0192 L10TWAXSH03 L2TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0193 L10TWAXSH03 L3TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0194 L10TWAXSH03 L4TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0195 L10TWAXSH03 L5TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0196 L10TWAXSH03 L6TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0197 L10TWAXSH03 L7TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0198 L10TWAXSH03 L8TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0199 L10TWAXSH03 L9TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0200 L10TWAXSH03 L10TWAXSH04 {max(min(M_stray002/sqrt(abs(LsS2_TWAXSH03*LsS2_TWAXSH04)),0.999),-0.999)}
Cstray002 CAPTWAXSH03 CAPTWAXSH04 {C_stray002} $ C#002=<C_stray002>
Kstray0201 L1TWAXSH01 L1TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)} $ M#003=<M_stray003>
Kstray0202 L1TWAXSH01 L2TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0203 L1TWAXSH01 L3TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0204 L1TWAXSH01 L4TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0205 L1TWAXSH01 L5TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0206 L1TWAXSH01 L6TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0207 L1TWAXSH01 L7TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0208 L1TWAXSH01 L8TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0209 L1TWAXSH01 L9TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0210 L1TWAXSH01 L10TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0211 L2TWAXSH01 L1TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0212 L2TWAXSH01 L2TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0213 L2TWAXSH01 L3TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0214 L2TWAXSH01 L4TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0215 L2TWAXSH01 L5TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0216 L2TWAXSH01 L6TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0217 L2TWAXSH01 L7TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0218 L2TWAXSH01 L8TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0219 L2TWAXSH01 L9TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0220 L2TWAXSH01 L10TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0221 L3TWAXSH01 L1TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0222 L3TWAXSH01 L2TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0223 L3TWAXSH01 L3TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0224 L3TWAXSH01 L4TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0225 L3TWAXSH01 L5TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0226 L3TWAXSH01 L6TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0227 L3TWAXSH01 L7TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0228 L3TWAXSH01 L8TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0229 L3TWAXSH01 L9TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0230 L3TWAXSH01 L10TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0231 L4TWAXSH01 L1TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0232 L4TWAXSH01 L2TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0233 L4TWAXSH01 L3TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0234 L4TWAXSH01 L4TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0235 L4TWAXSH01 L5TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0236 L4TWAXSH01 L6TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0237 L4TWAXSH01 L7TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0238 L4TWAXSH01 L8TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0239 L4TWAXSH01 L9TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0240 L4TWAXSH01 L10TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0241 L5TWAXSH01 L1TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0242 L5TWAXSH01 L2TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0243 L5TWAXSH01 L3TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0244 L5TWAXSH01 L4TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0245 L5TWAXSH01 L5TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0246 L5TWAXSH01 L6TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0247 L5TWAXSH01 L7TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0248 L5TWAXSH01 L8TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0249 L5TWAXSH01 L9TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0250 L5TWAXSH01 L10TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0251 L6TWAXSH01 L1TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0252 L6TWAXSH01 L2TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0253 L6TWAXSH01 L3TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0254 L6TWAXSH01 L4TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0255 L6TWAXSH01 L5TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0256 L6TWAXSH01 L6TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0257 L6TWAXSH01 L7TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0258 L6TWAXSH01 L8TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0259 L6TWAXSH01 L9TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0260 L6TWAXSH01 L10TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0261 L7TWAXSH01 L1TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0262 L7TWAXSH01 L2TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0263 L7TWAXSH01 L3TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0264 L7TWAXSH01 L4TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0265 L7TWAXSH01 L5TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0266 L7TWAXSH01 L6TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0267 L7TWAXSH01 L7TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0268 L7TWAXSH01 L8TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0269 L7TWAXSH01 L9TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0270 L7TWAXSH01 L10TWAXSH03 {max(min(M_stray003/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0271 L8TWAXSH01 L1TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0272 L8TWAXSH01 L2TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0273 L8TWAXSH01 L3TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0274 L8TWAXSH01 L4TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0275 L8TWAXSH01 L5TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0276 L8TWAXSH01 L6TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0277 L8TWAXSH01 L7TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0278 L8TWAXSH01 L8TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0279 L8TWAXSH01 L9TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0280 L8TWAXSH01 L10TWAXSH03 {max(min(M_stray003/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0281 L9TWAXSH01 L1TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0282 L9TWAXSH01 L2TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0283 L9TWAXSH01 L3TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0284 L9TWAXSH01 L4TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0285 L9TWAXSH01 L5TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0286 L9TWAXSH01 L6TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0287 L9TWAXSH01 L7TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0288 L9TWAXSH01 L8TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0289 L9TWAXSH01 L9TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0290 L9TWAXSH01 L10TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0291 L10TWAXSH01 L1TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0292 L10TWAXSH01 L2TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0293 L10TWAXSH01 L3TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0294 L10TWAXSH01 L4TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0295 L10TWAXSH01 L5TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0296 L10TWAXSH01 L6TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0297 L10TWAXSH01 L7TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0298 L10TWAXSH01 L8TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0299 L10TWAXSH01 L9TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0300 L10TWAXSH01 L10TWAXSH03 {max(min(M_stray003/sqrt(abs(LsS2_TWAXSH01*LsS2_TWAXSH03)),0.999),-0.999)}
Cstray003 CAPTWAXSH01 CAPTWAXSH03 {C_stray003} $ C#003=<C_stray003>
Kstray0301 L1TWAXSH01 L1TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)} $ M#003=<M_stray004>
Kstray0302 L1TWAXSH01 L2TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0303 L1TWAXSH01 L3TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0304 L1TWAXSH01 L4TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0305 L1TWAXSH01 L5TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0306 L1TWAXSH01 L6TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0307 L1TWAXSH01 L7TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0308 L1TWAXSH01 L8TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0309 L1TWAXSH01 L9TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0310 L1TWAXSH01 L10TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0311 L2TWAXSH01 L1TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0312 L2TWAXSH01 L2TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0313 L2TWAXSH01 L3TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0314 L2TWAXSH01 L4TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0315 L2TWAXSH01 L5TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0316 L2TWAXSH01 L6TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0317 L2TWAXSH01 L7TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0318 L2TWAXSH01 L8TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0319 L2TWAXSH01 L9TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0320 L2TWAXSH01 L10TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0321 L3TWAXSH01 L1TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0322 L3TWAXSH01 L2TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0323 L3TWAXSH01 L3TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0324 L3TWAXSH01 L4TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0325 L3TWAXSH01 L5TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0326 L3TWAXSH01 L6TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0327 L3TWAXSH01 L7TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0328 L3TWAXSH01 L8TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0329 L3TWAXSH01 L9TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0330 L3TWAXSH01 L10TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0331 L4TWAXSH01 L1TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0332 L4TWAXSH01 L2TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0333 L4TWAXSH01 L3TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0334 L4TWAXSH01 L4TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0335 L4TWAXSH01 L5TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0336 L4TWAXSH01 L6TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0337 L4TWAXSH01 L7TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0338 L4TWAXSH01 L8TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0339 L4TWAXSH01 L9TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0340 L4TWAXSH01 L10TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0341 L5TWAXSH01 L1TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0342 L5TWAXSH01 L2TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0343 L5TWAXSH01 L3TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0344 L5TWAXSH01 L4TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0345 L5TWAXSH01 L5TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0346 L5TWAXSH01 L6TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0347 L5TWAXSH01 L7TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0348 L5TWAXSH01 L8TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0349 L5TWAXSH01 L9TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0350 L5TWAXSH01 L10TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0351 L6TWAXSH01 L1TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0352 L6TWAXSH01 L2TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0353 L6TWAXSH01 L3TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0354 L6TWAXSH01 L4TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0355 L6TWAXSH01 L5TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0356 L6TWAXSH01 L6TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0357 L6TWAXSH01 L7TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0358 L6TWAXSH01 L8TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0359 L6TWAXSH01 L9TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0360 L6TWAXSH01 L10TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0361 L7TWAXSH01 L1TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0362 L7TWAXSH01 L2TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0363 L7TWAXSH01 L3TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0364 L7TWAXSH01 L4TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0365 L7TWAXSH01 L5TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0366 L7TWAXSH01 L6TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0367 L7TWAXSH01 L7TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0368 L7TWAXSH01 L8TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0369 L7TWAXSH01 L9TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0370 L7TWAXSH01 L10TWAXSH04 {max(min(M_stray004/sqrt(abs(Ls2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0371 L8TWAXSH01 L1TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0372 L8TWAXSH01 L2TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0373 L8TWAXSH01 L3TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0374 L8TWAXSH01 L4TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0375 L8TWAXSH01 L5TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0376 L8TWAXSH01 L6TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0377 L8TWAXSH01 L7TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0378 L8TWAXSH01 L8TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0379 L8TWAXSH01 L9TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0380 L8TWAXSH01 L10TWAXSH04 {max(min(M_stray004/sqrt(abs(LsG2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0381 L9TWAXSH01 L1TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0382 L9TWAXSH01 L2TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0383 L9TWAXSH01 L3TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0384 L9TWAXSH01 L4TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0385 L9TWAXSH01 L5TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0386 L9TWAXSH01 L6TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0387 L9TWAXSH01 L7TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0388 L9TWAXSH01 L8TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0389 L9TWAXSH01 L9TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0390 L9TWAXSH01 L10TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0391 L10TWAXSH01 L1TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0392 L10TWAXSH01 L2TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0393 L10TWAXSH01 L3TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0394 L10TWAXSH01 L4TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0395 L10TWAXSH01 L5TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0396 L10TWAXSH01 L6TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0397 L10TWAXSH01 L7TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0398 L10TWAXSH01 L8TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0399 L10TWAXSH01 L9TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0400 L10TWAXSH01 L10TWAXSH04 {max(min(M_stray004/sqrt(abs(LsS2_TWAXSH01*LsS2_TWAXSH04)),0.999),-0.999)}
Cstray004 CAPTWAXSH01 CAPTWAXSH04 {C_stray004} $ C#003=<C_stray004>
Kstray0401 L1TWAXSH02 L1TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)} $ M#003=<M_stray005>
Kstray0402 L1TWAXSH02 L2TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0403 L1TWAXSH02 L3TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0404 L1TWAXSH02 L4TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0405 L1TWAXSH02 L5TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0406 L1TWAXSH02 L6TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0407 L1TWAXSH02 L7TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0408 L1TWAXSH02 L8TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0409 L1TWAXSH02 L9TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0410 L1TWAXSH02 L10TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0411 L2TWAXSH02 L1TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0412 L2TWAXSH02 L2TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0413 L2TWAXSH02 L3TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0414 L2TWAXSH02 L4TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0415 L2TWAXSH02 L5TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0416 L2TWAXSH02 L6TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0417 L2TWAXSH02 L7TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0418 L2TWAXSH02 L8TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0419 L2TWAXSH02 L9TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0420 L2TWAXSH02 L10TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0421 L3TWAXSH02 L1TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0422 L3TWAXSH02 L2TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0423 L3TWAXSH02 L3TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0424 L3TWAXSH02 L4TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0425 L3TWAXSH02 L5TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0426 L3TWAXSH02 L6TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0427 L3TWAXSH02 L7TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0428 L3TWAXSH02 L8TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0429 L3TWAXSH02 L9TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0430 L3TWAXSH02 L10TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0431 L4TWAXSH02 L1TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0432 L4TWAXSH02 L2TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0433 L4TWAXSH02 L3TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0434 L4TWAXSH02 L4TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0435 L4TWAXSH02 L5TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0436 L4TWAXSH02 L6TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0437 L4TWAXSH02 L7TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0438 L4TWAXSH02 L8TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0439 L4TWAXSH02 L9TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0440 L4TWAXSH02 L10TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0441 L5TWAXSH02 L1TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0442 L5TWAXSH02 L2TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0443 L5TWAXSH02 L3TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0444 L5TWAXSH02 L4TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0445 L5TWAXSH02 L5TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0446 L5TWAXSH02 L6TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0447 L5TWAXSH02 L7TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0448 L5TWAXSH02 L8TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0449 L5TWAXSH02 L9TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0450 L5TWAXSH02 L10TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0451 L6TWAXSH02 L1TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0452 L6TWAXSH02 L2TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0453 L6TWAXSH02 L3TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0454 L6TWAXSH02 L4TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0455 L6TWAXSH02 L5TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0456 L6TWAXSH02 L6TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0457 L6TWAXSH02 L7TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0458 L6TWAXSH02 L8TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0459 L6TWAXSH02 L9TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0460 L6TWAXSH02 L10TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0461 L7TWAXSH02 L1TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0462 L7TWAXSH02 L2TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0463 L7TWAXSH02 L3TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0464 L7TWAXSH02 L4TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0465 L7TWAXSH02 L5TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0466 L7TWAXSH02 L6TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0467 L7TWAXSH02 L7TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0468 L7TWAXSH02 L8TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0469 L7TWAXSH02 L9TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0470 L7TWAXSH02 L10TWAXSH03 {max(min(M_stray005/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0471 L8TWAXSH02 L1TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0472 L8TWAXSH02 L2TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0473 L8TWAXSH02 L3TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0474 L8TWAXSH02 L4TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0475 L8TWAXSH02 L5TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0476 L8TWAXSH02 L6TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0477 L8TWAXSH02 L7TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0478 L8TWAXSH02 L8TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0479 L8TWAXSH02 L9TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0480 L8TWAXSH02 L10TWAXSH03 {max(min(M_stray005/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0481 L9TWAXSH02 L1TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0482 L9TWAXSH02 L2TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0483 L9TWAXSH02 L3TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0484 L9TWAXSH02 L4TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0485 L9TWAXSH02 L5TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0486 L9TWAXSH02 L6TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0487 L9TWAXSH02 L7TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0488 L9TWAXSH02 L8TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0489 L9TWAXSH02 L9TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0490 L9TWAXSH02 L10TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0491 L10TWAXSH02 L1TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0492 L10TWAXSH02 L2TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0493 L10TWAXSH02 L3TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0494 L10TWAXSH02 L4TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0495 L10TWAXSH02 L5TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0496 L10TWAXSH02 L6TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0497 L10TWAXSH02 L7TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray0498 L10TWAXSH02 L8TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray0499 L10TWAXSH02 L9TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray0500 L10TWAXSH02 L10TWAXSH03 {max(min(M_stray005/sqrt(abs(LsS2_TWAXSH02*LsS2_TWAXSH03)),0.999),-0.999)}
Cstray005 CAPTWAXSH02 CAPTWAXSH03 {C_stray005} $ C#003=<C_stray005>
Kstray0501 L1TWAXSH02 L1TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)} $ M#003=<M_stray006>
Kstray0502 L1TWAXSH02 L2TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0503 L1TWAXSH02 L3TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0504 L1TWAXSH02 L4TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0505 L1TWAXSH02 L5TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0506 L1TWAXSH02 L6TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0507 L1TWAXSH02 L7TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0508 L1TWAXSH02 L8TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0509 L1TWAXSH02 L9TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0510 L1TWAXSH02 L10TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0511 L2TWAXSH02 L1TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0512 L2TWAXSH02 L2TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0513 L2TWAXSH02 L3TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0514 L2TWAXSH02 L4TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0515 L2TWAXSH02 L5TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0516 L2TWAXSH02 L6TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0517 L2TWAXSH02 L7TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0518 L2TWAXSH02 L8TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0519 L2TWAXSH02 L9TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0520 L2TWAXSH02 L10TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0521 L3TWAXSH02 L1TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0522 L3TWAXSH02 L2TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0523 L3TWAXSH02 L3TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0524 L3TWAXSH02 L4TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0525 L3TWAXSH02 L5TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0526 L3TWAXSH02 L6TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0527 L3TWAXSH02 L7TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0528 L3TWAXSH02 L8TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0529 L3TWAXSH02 L9TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0530 L3TWAXSH02 L10TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0531 L4TWAXSH02 L1TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0532 L4TWAXSH02 L2TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0533 L4TWAXSH02 L3TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0534 L4TWAXSH02 L4TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0535 L4TWAXSH02 L5TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0536 L4TWAXSH02 L6TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0537 L4TWAXSH02 L7TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0538 L4TWAXSH02 L8TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0539 L4TWAXSH02 L9TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0540 L4TWAXSH02 L10TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0541 L5TWAXSH02 L1TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0542 L5TWAXSH02 L2TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0543 L5TWAXSH02 L3TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0544 L5TWAXSH02 L4TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0545 L5TWAXSH02 L5TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0546 L5TWAXSH02 L6TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0547 L5TWAXSH02 L7TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0548 L5TWAXSH02 L8TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0549 L5TWAXSH02 L9TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0550 L5TWAXSH02 L10TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0551 L6TWAXSH02 L1TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0552 L6TWAXSH02 L2TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0553 L6TWAXSH02 L3TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0554 L6TWAXSH02 L4TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0555 L6TWAXSH02 L5TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0556 L6TWAXSH02 L6TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0557 L6TWAXSH02 L7TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0558 L6TWAXSH02 L8TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0559 L6TWAXSH02 L9TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0560 L6TWAXSH02 L10TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0561 L7TWAXSH02 L1TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0562 L7TWAXSH02 L2TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0563 L7TWAXSH02 L3TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0564 L7TWAXSH02 L4TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0565 L7TWAXSH02 L5TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0566 L7TWAXSH02 L6TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0567 L7TWAXSH02 L7TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0568 L7TWAXSH02 L8TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0569 L7TWAXSH02 L9TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0570 L7TWAXSH02 L10TWAXSH04 {max(min(M_stray006/sqrt(abs(Ls2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0571 L8TWAXSH02 L1TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0572 L8TWAXSH02 L2TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0573 L8TWAXSH02 L3TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0574 L8TWAXSH02 L4TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0575 L8TWAXSH02 L5TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0576 L8TWAXSH02 L6TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0577 L8TWAXSH02 L7TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0578 L8TWAXSH02 L8TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0579 L8TWAXSH02 L9TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0580 L8TWAXSH02 L10TWAXSH04 {max(min(M_stray006/sqrt(abs(LsG2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0581 L9TWAXSH02 L1TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0582 L9TWAXSH02 L2TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0583 L9TWAXSH02 L3TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0584 L9TWAXSH02 L4TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0585 L9TWAXSH02 L5TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0586 L9TWAXSH02 L6TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0587 L9TWAXSH02 L7TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0588 L9TWAXSH02 L8TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0589 L9TWAXSH02 L9TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0590 L9TWAXSH02 L10TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0591 L10TWAXSH02 L1TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0592 L10TWAXSH02 L2TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0593 L10TWAXSH02 L3TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0594 L10TWAXSH02 L4TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0595 L10TWAXSH02 L5TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0596 L10TWAXSH02 L6TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0597 L10TWAXSH02 L7TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray0598 L10TWAXSH02 L8TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray0599 L10TWAXSH02 L9TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray0600 L10TWAXSH02 L10TWAXSH04 {max(min(M_stray006/sqrt(abs(LsS2_TWAXSH02*LsS2_TWAXSH04)),0.999),-0.999)}
Cstray006 CAPTWAXSH02 CAPTWAXSH04 {C_stray006} $ C#003=<C_stray006>
Kstray0601 L1TWAXSH01 L1COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)} $ M#004=<M_stray007>
Kstray0602 L1TWAXSH01 L2COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0603 L1TWAXSH01 L3COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0604 L1TWAXSH01 L4COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0605 L2TWAXSH01 L1COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0606 L2TWAXSH01 L2COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0607 L2TWAXSH01 L3COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0608 L2TWAXSH01 L4COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0609 L3TWAXSH01 L1COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0610 L3TWAXSH01 L2COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0611 L3TWAXSH01 L3COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0612 L3TWAXSH01 L4COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0613 L4TWAXSH01 L1COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0614 L4TWAXSH01 L2COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0615 L4TWAXSH01 L3COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0616 L4TWAXSH01 L4COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0617 L5TWAXSH01 L1COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0618 L5TWAXSH01 L2COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0619 L5TWAXSH01 L3COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0620 L5TWAXSH01 L4COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0621 L6TWAXSH01 L1COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0622 L6TWAXSH01 L2COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0623 L6TWAXSH01 L3COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0624 L6TWAXSH01 L4COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0625 L7TWAXSH01 L1COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0626 L7TWAXSH01 L2COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0627 L7TWAXSH01 L3COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0628 L7TWAXSH01 L4COAXCAB03 {max(min(M_stray007/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0629 L8TWAXSH01 L1COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0630 L8TWAXSH01 L2COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0631 L8TWAXSH01 L3COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0632 L8TWAXSH01 L4COAXCAB03 {max(min(M_stray007/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0633 L9TWAXSH01 L1COAXCAB03 {max(min(M_stray007/sqrt(abs(LsS2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0634 L9TWAXSH01 L2COAXCAB03 {max(min(M_stray007/sqrt(abs(LsS2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0635 L9TWAXSH01 L3COAXCAB03 {max(min(M_stray007/sqrt(abs(LsS2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0636 L9TWAXSH01 L4COAXCAB03 {max(min(M_stray007/sqrt(abs(LsS2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0637 L10TWAXSH01 L1COAXCAB03 {max(min(M_stray007/sqrt(abs(LsS2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0638 L10TWAXSH01 L2COAXCAB03 {max(min(M_stray007/sqrt(abs(LsS2_TWAXSH01*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0639 L10TWAXSH01 L3COAXCAB03 {max(min(M_stray007/sqrt(abs(LsS2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0640 L10TWAXSH01 L4COAXCAB03 {max(min(M_stray007/sqrt(abs(LsS2_TWAXSH01*LsG2_COAXCAB03)),0.999),-0.999)}
Cstray007 CAPTWAXSH01 n005COAXCAB03 {C_stray007} $ C#004=<C_stray007>
Kstray0641 L1TWAXSH02 L1COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)} $ M#004=<M_stray008>
Kstray0642 L1TWAXSH02 L2COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0643 L1TWAXSH02 L3COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0644 L1TWAXSH02 L4COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0645 L2TWAXSH02 L1COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0646 L2TWAXSH02 L2COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0647 L2TWAXSH02 L3COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0648 L2TWAXSH02 L4COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0649 L3TWAXSH02 L1COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0650 L3TWAXSH02 L2COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0651 L3TWAXSH02 L3COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0652 L3TWAXSH02 L4COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0653 L4TWAXSH02 L1COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0654 L4TWAXSH02 L2COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0655 L4TWAXSH02 L3COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0656 L4TWAXSH02 L4COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0657 L5TWAXSH02 L1COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0658 L5TWAXSH02 L2COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0659 L5TWAXSH02 L3COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0660 L5TWAXSH02 L4COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0661 L6TWAXSH02 L1COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0662 L6TWAXSH02 L2COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0663 L6TWAXSH02 L3COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0664 L6TWAXSH02 L4COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0665 L7TWAXSH02 L1COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0666 L7TWAXSH02 L2COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0667 L7TWAXSH02 L3COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0668 L7TWAXSH02 L4COAXCAB03 {max(min(M_stray008/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0669 L8TWAXSH02 L1COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0670 L8TWAXSH02 L2COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0671 L8TWAXSH02 L3COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0672 L8TWAXSH02 L4COAXCAB03 {max(min(M_stray008/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0673 L9TWAXSH02 L1COAXCAB03 {max(min(M_stray008/sqrt(abs(LsS2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0674 L9TWAXSH02 L2COAXCAB03 {max(min(M_stray008/sqrt(abs(LsS2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0675 L9TWAXSH02 L3COAXCAB03 {max(min(M_stray008/sqrt(abs(LsS2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0676 L9TWAXSH02 L4COAXCAB03 {max(min(M_stray008/sqrt(abs(LsS2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0677 L10TWAXSH02 L1COAXCAB03 {max(min(M_stray008/sqrt(abs(LsS2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0678 L10TWAXSH02 L2COAXCAB03 {max(min(M_stray008/sqrt(abs(LsS2_TWAXSH02*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0679 L10TWAXSH02 L3COAXCAB03 {max(min(M_stray008/sqrt(abs(LsS2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0680 L10TWAXSH02 L4COAXCAB03 {max(min(M_stray008/sqrt(abs(LsS2_TWAXSH02*LsG2_COAXCAB03)),0.999),-0.999)}
Cstray008 CAPTWAXSH02 n005COAXCAB03 {C_stray008} $ C#004=<C_stray008>
Kstray0681 L1TWAXSH03 L1COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)} $ M#004=<M_stray009>
Kstray0682 L1TWAXSH03 L2COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0683 L1TWAXSH03 L3COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0684 L1TWAXSH03 L4COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0685 L2TWAXSH03 L1COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0686 L2TWAXSH03 L2COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0687 L2TWAXSH03 L3COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0688 L2TWAXSH03 L4COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0689 L3TWAXSH03 L1COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0690 L3TWAXSH03 L2COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0691 L3TWAXSH03 L3COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0692 L3TWAXSH03 L4COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0693 L4TWAXSH03 L1COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0694 L4TWAXSH03 L2COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0695 L4TWAXSH03 L3COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0696 L4TWAXSH03 L4COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0697 L5TWAXSH03 L1COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0698 L5TWAXSH03 L2COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0699 L5TWAXSH03 L3COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0700 L5TWAXSH03 L4COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0701 L6TWAXSH03 L1COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0702 L6TWAXSH03 L2COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0703 L6TWAXSH03 L3COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0704 L6TWAXSH03 L4COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0705 L7TWAXSH03 L1COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0706 L7TWAXSH03 L2COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0707 L7TWAXSH03 L3COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0708 L7TWAXSH03 L4COAXCAB03 {max(min(M_stray009/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0709 L8TWAXSH03 L1COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0710 L8TWAXSH03 L2COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0711 L8TWAXSH03 L3COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0712 L8TWAXSH03 L4COAXCAB03 {max(min(M_stray009/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0713 L9TWAXSH03 L1COAXCAB03 {max(min(M_stray009/sqrt(abs(LsS2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0714 L9TWAXSH03 L2COAXCAB03 {max(min(M_stray009/sqrt(abs(LsS2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0715 L9TWAXSH03 L3COAXCAB03 {max(min(M_stray009/sqrt(abs(LsS2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0716 L9TWAXSH03 L4COAXCAB03 {max(min(M_stray009/sqrt(abs(LsS2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0717 L10TWAXSH03 L1COAXCAB03 {max(min(M_stray009/sqrt(abs(LsS2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0718 L10TWAXSH03 L2COAXCAB03 {max(min(M_stray009/sqrt(abs(LsS2_TWAXSH03*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0719 L10TWAXSH03 L3COAXCAB03 {max(min(M_stray009/sqrt(abs(LsS2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0720 L10TWAXSH03 L4COAXCAB03 {max(min(M_stray009/sqrt(abs(LsS2_TWAXSH03*LsG2_COAXCAB03)),0.999),-0.999)}
Cstray009 CAPTWAXSH03 n005COAXCAB03 {C_stray009} $ C#004=<C_stray009>
Kstray0721 L1TWAXSH04 L1COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)} $ M#004=<M_stray010>
Kstray0722 L1TWAXSH04 L2COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0723 L1TWAXSH04 L3COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0724 L1TWAXSH04 L4COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0725 L2TWAXSH04 L1COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0726 L2TWAXSH04 L2COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0727 L2TWAXSH04 L3COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0728 L2TWAXSH04 L4COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0729 L3TWAXSH04 L1COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0730 L3TWAXSH04 L2COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0731 L3TWAXSH04 L3COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0732 L3TWAXSH04 L4COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0733 L4TWAXSH04 L1COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0734 L4TWAXSH04 L2COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0735 L4TWAXSH04 L3COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0736 L4TWAXSH04 L4COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0737 L5TWAXSH04 L1COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0738 L5TWAXSH04 L2COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0739 L5TWAXSH04 L3COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0740 L5TWAXSH04 L4COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0741 L6TWAXSH04 L1COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0742 L6TWAXSH04 L2COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0743 L6TWAXSH04 L3COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0744 L6TWAXSH04 L4COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0745 L7TWAXSH04 L1COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0746 L7TWAXSH04 L2COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0747 L7TWAXSH04 L3COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0748 L7TWAXSH04 L4COAXCAB03 {max(min(M_stray010/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0749 L8TWAXSH04 L1COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0750 L8TWAXSH04 L2COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0751 L8TWAXSH04 L3COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0752 L8TWAXSH04 L4COAXCAB03 {max(min(M_stray010/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0753 L9TWAXSH04 L1COAXCAB03 {max(min(M_stray010/sqrt(abs(LsS2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0754 L9TWAXSH04 L2COAXCAB03 {max(min(M_stray010/sqrt(abs(LsS2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0755 L9TWAXSH04 L3COAXCAB03 {max(min(M_stray010/sqrt(abs(LsS2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0756 L9TWAXSH04 L4COAXCAB03 {max(min(M_stray010/sqrt(abs(LsS2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0757 L10TWAXSH04 L1COAXCAB03 {max(min(M_stray010/sqrt(abs(LsS2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0758 L10TWAXSH04 L2COAXCAB03 {max(min(M_stray010/sqrt(abs(LsS2_TWAXSH04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray0759 L10TWAXSH04 L3COAXCAB03 {max(min(M_stray010/sqrt(abs(LsS2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray0760 L10TWAXSH04 L4COAXCAB03 {max(min(M_stray010/sqrt(abs(LsS2_TWAXSH04*LsG2_COAXCAB03)),0.999),-0.999)}
Cstray010 CAPTWAXSH04 n005COAXCAB03 {C_stray010} $ C#004=<C_stray010>
Kstray0761 L1TWAXSH01 L1COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)} $ M#005=<M_stray011>
Kstray0762 L1TWAXSH01 L2COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0763 L1TWAXSH01 L3COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0764 L1TWAXSH01 L4COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0765 L2TWAXSH01 L1COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0766 L2TWAXSH01 L2COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0767 L2TWAXSH01 L3COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0768 L2TWAXSH01 L4COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0769 L3TWAXSH01 L1COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0770 L3TWAXSH01 L2COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0771 L3TWAXSH01 L3COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0772 L3TWAXSH01 L4COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0773 L4TWAXSH01 L1COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0774 L4TWAXSH01 L2COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0775 L4TWAXSH01 L3COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0776 L4TWAXSH01 L4COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0777 L5TWAXSH01 L1COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0778 L5TWAXSH01 L2COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0779 L5TWAXSH01 L3COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0780 L5TWAXSH01 L4COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0781 L6TWAXSH01 L1COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0782 L6TWAXSH01 L2COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0783 L6TWAXSH01 L3COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0784 L6TWAXSH01 L4COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0785 L7TWAXSH01 L1COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0786 L7TWAXSH01 L2COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0787 L7TWAXSH01 L3COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0788 L7TWAXSH01 L4COAXCAB02 {max(min(M_stray011/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0789 L8TWAXSH01 L1COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0790 L8TWAXSH01 L2COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0791 L8TWAXSH01 L3COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0792 L8TWAXSH01 L4COAXCAB02 {max(min(M_stray011/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0793 L9TWAXSH01 L1COAXCAB02 {max(min(M_stray011/sqrt(abs(LsS2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0794 L9TWAXSH01 L2COAXCAB02 {max(min(M_stray011/sqrt(abs(LsS2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0795 L9TWAXSH01 L3COAXCAB02 {max(min(M_stray011/sqrt(abs(LsS2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0796 L9TWAXSH01 L4COAXCAB02 {max(min(M_stray011/sqrt(abs(LsS2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0797 L10TWAXSH01 L1COAXCAB02 {max(min(M_stray011/sqrt(abs(LsS2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0798 L10TWAXSH01 L2COAXCAB02 {max(min(M_stray011/sqrt(abs(LsS2_TWAXSH01*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0799 L10TWAXSH01 L3COAXCAB02 {max(min(M_stray011/sqrt(abs(LsS2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0800 L10TWAXSH01 L4COAXCAB02 {max(min(M_stray011/sqrt(abs(LsS2_TWAXSH01*LsG2_COAXCAB02)),0.999),-0.999)}
Cstray011 CAPTWAXSH01 n005COAXCAB02 {C_stray011} $ C#005=<C_stray011>
Kstray0801 L1TWAXSH01 L1COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)} $ M#005=<M_stray012>
Kstray0802 L1TWAXSH01 L2COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0803 L1TWAXSH01 L3COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0804 L1TWAXSH01 L4COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0805 L2TWAXSH01 L1COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0806 L2TWAXSH01 L2COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0807 L2TWAXSH01 L3COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0808 L2TWAXSH01 L4COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0809 L3TWAXSH01 L1COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0810 L3TWAXSH01 L2COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0811 L3TWAXSH01 L3COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0812 L3TWAXSH01 L4COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0813 L4TWAXSH01 L1COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0814 L4TWAXSH01 L2COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0815 L4TWAXSH01 L3COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0816 L4TWAXSH01 L4COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0817 L5TWAXSH01 L1COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0818 L5TWAXSH01 L2COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0819 L5TWAXSH01 L3COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0820 L5TWAXSH01 L4COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0821 L6TWAXSH01 L1COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0822 L6TWAXSH01 L2COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0823 L6TWAXSH01 L3COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0824 L6TWAXSH01 L4COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0825 L7TWAXSH01 L1COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0826 L7TWAXSH01 L2COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0827 L7TWAXSH01 L3COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0828 L7TWAXSH01 L4COAXCAB01 {max(min(M_stray012/sqrt(abs(Ls2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0829 L8TWAXSH01 L1COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0830 L8TWAXSH01 L2COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0831 L8TWAXSH01 L3COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0832 L8TWAXSH01 L4COAXCAB01 {max(min(M_stray012/sqrt(abs(LsG2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0833 L9TWAXSH01 L1COAXCAB01 {max(min(M_stray012/sqrt(abs(LsS2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0834 L9TWAXSH01 L2COAXCAB01 {max(min(M_stray012/sqrt(abs(LsS2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0835 L9TWAXSH01 L3COAXCAB01 {max(min(M_stray012/sqrt(abs(LsS2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0836 L9TWAXSH01 L4COAXCAB01 {max(min(M_stray012/sqrt(abs(LsS2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0837 L10TWAXSH01 L1COAXCAB01 {max(min(M_stray012/sqrt(abs(LsS2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0838 L10TWAXSH01 L2COAXCAB01 {max(min(M_stray012/sqrt(abs(LsS2_TWAXSH01*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0839 L10TWAXSH01 L3COAXCAB01 {max(min(M_stray012/sqrt(abs(LsS2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0840 L10TWAXSH01 L4COAXCAB01 {max(min(M_stray012/sqrt(abs(LsS2_TWAXSH01*LsG2_COAXCAB01)),0.999),-0.999)}
Cstray012 CAPTWAXSH01 n005COAXCAB01 {C_stray012} $ C#005=<C_stray012>
Kstray0841 L1TWAXSH02 L1COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)} $ M#005=<M_stray013>
Kstray0842 L1TWAXSH02 L2COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0843 L1TWAXSH02 L3COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0844 L1TWAXSH02 L4COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0845 L2TWAXSH02 L1COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0846 L2TWAXSH02 L2COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0847 L2TWAXSH02 L3COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0848 L2TWAXSH02 L4COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0849 L3TWAXSH02 L1COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0850 L3TWAXSH02 L2COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0851 L3TWAXSH02 L3COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0852 L3TWAXSH02 L4COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0853 L4TWAXSH02 L1COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0854 L4TWAXSH02 L2COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0855 L4TWAXSH02 L3COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0856 L4TWAXSH02 L4COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0857 L5TWAXSH02 L1COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0858 L5TWAXSH02 L2COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0859 L5TWAXSH02 L3COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0860 L5TWAXSH02 L4COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0861 L6TWAXSH02 L1COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0862 L6TWAXSH02 L2COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0863 L6TWAXSH02 L3COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0864 L6TWAXSH02 L4COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0865 L7TWAXSH02 L1COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0866 L7TWAXSH02 L2COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0867 L7TWAXSH02 L3COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0868 L7TWAXSH02 L4COAXCAB02 {max(min(M_stray013/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0869 L8TWAXSH02 L1COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0870 L8TWAXSH02 L2COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0871 L8TWAXSH02 L3COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0872 L8TWAXSH02 L4COAXCAB02 {max(min(M_stray013/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0873 L9TWAXSH02 L1COAXCAB02 {max(min(M_stray013/sqrt(abs(LsS2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0874 L9TWAXSH02 L2COAXCAB02 {max(min(M_stray013/sqrt(abs(LsS2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0875 L9TWAXSH02 L3COAXCAB02 {max(min(M_stray013/sqrt(abs(LsS2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0876 L9TWAXSH02 L4COAXCAB02 {max(min(M_stray013/sqrt(abs(LsS2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0877 L10TWAXSH02 L1COAXCAB02 {max(min(M_stray013/sqrt(abs(LsS2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0878 L10TWAXSH02 L2COAXCAB02 {max(min(M_stray013/sqrt(abs(LsS2_TWAXSH02*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0879 L10TWAXSH02 L3COAXCAB02 {max(min(M_stray013/sqrt(abs(LsS2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0880 L10TWAXSH02 L4COAXCAB02 {max(min(M_stray013/sqrt(abs(LsS2_TWAXSH02*LsG2_COAXCAB02)),0.999),-0.999)}
Cstray013 CAPTWAXSH02 n005COAXCAB02 {C_stray013} $ C#005=<C_stray013>
Kstray0881 L1TWAXSH02 L1COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)} $ M#005=<M_stray014>
Kstray0882 L1TWAXSH02 L2COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0883 L1TWAXSH02 L3COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0884 L1TWAXSH02 L4COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0885 L2TWAXSH02 L1COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0886 L2TWAXSH02 L2COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0887 L2TWAXSH02 L3COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0888 L2TWAXSH02 L4COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0889 L3TWAXSH02 L1COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0890 L3TWAXSH02 L2COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0891 L3TWAXSH02 L3COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0892 L3TWAXSH02 L4COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0893 L4TWAXSH02 L1COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0894 L4TWAXSH02 L2COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0895 L4TWAXSH02 L3COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0896 L4TWAXSH02 L4COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0897 L5TWAXSH02 L1COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0898 L5TWAXSH02 L2COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0899 L5TWAXSH02 L3COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0900 L5TWAXSH02 L4COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0901 L6TWAXSH02 L1COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0902 L6TWAXSH02 L2COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0903 L6TWAXSH02 L3COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0904 L6TWAXSH02 L4COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0905 L7TWAXSH02 L1COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0906 L7TWAXSH02 L2COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0907 L7TWAXSH02 L3COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0908 L7TWAXSH02 L4COAXCAB01 {max(min(M_stray014/sqrt(abs(Ls2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0909 L8TWAXSH02 L1COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0910 L8TWAXSH02 L2COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0911 L8TWAXSH02 L3COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0912 L8TWAXSH02 L4COAXCAB01 {max(min(M_stray014/sqrt(abs(LsG2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0913 L9TWAXSH02 L1COAXCAB01 {max(min(M_stray014/sqrt(abs(LsS2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0914 L9TWAXSH02 L2COAXCAB01 {max(min(M_stray014/sqrt(abs(LsS2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0915 L9TWAXSH02 L3COAXCAB01 {max(min(M_stray014/sqrt(abs(LsS2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0916 L9TWAXSH02 L4COAXCAB01 {max(min(M_stray014/sqrt(abs(LsS2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0917 L10TWAXSH02 L1COAXCAB01 {max(min(M_stray014/sqrt(abs(LsS2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0918 L10TWAXSH02 L2COAXCAB01 {max(min(M_stray014/sqrt(abs(LsS2_TWAXSH02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0919 L10TWAXSH02 L3COAXCAB01 {max(min(M_stray014/sqrt(abs(LsS2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0920 L10TWAXSH02 L4COAXCAB01 {max(min(M_stray014/sqrt(abs(LsS2_TWAXSH02*LsG2_COAXCAB01)),0.999),-0.999)}
Cstray014 CAPTWAXSH02 n005COAXCAB01 {C_stray014} $ C#005=<C_stray014>
Kstray0921 L1TWAXSH03 L1COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)} $ M#005=<M_stray015>
Kstray0922 L1TWAXSH03 L2COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0923 L1TWAXSH03 L3COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0924 L1TWAXSH03 L4COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0925 L2TWAXSH03 L1COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0926 L2TWAXSH03 L2COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0927 L2TWAXSH03 L3COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0928 L2TWAXSH03 L4COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0929 L3TWAXSH03 L1COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0930 L3TWAXSH03 L2COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0931 L3TWAXSH03 L3COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0932 L3TWAXSH03 L4COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0933 L4TWAXSH03 L1COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0934 L4TWAXSH03 L2COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0935 L4TWAXSH03 L3COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0936 L4TWAXSH03 L4COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0937 L5TWAXSH03 L1COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0938 L5TWAXSH03 L2COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0939 L5TWAXSH03 L3COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0940 L5TWAXSH03 L4COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0941 L6TWAXSH03 L1COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0942 L6TWAXSH03 L2COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0943 L6TWAXSH03 L3COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0944 L6TWAXSH03 L4COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0945 L7TWAXSH03 L1COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0946 L7TWAXSH03 L2COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0947 L7TWAXSH03 L3COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0948 L7TWAXSH03 L4COAXCAB02 {max(min(M_stray015/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0949 L8TWAXSH03 L1COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0950 L8TWAXSH03 L2COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0951 L8TWAXSH03 L3COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0952 L8TWAXSH03 L4COAXCAB02 {max(min(M_stray015/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0953 L9TWAXSH03 L1COAXCAB02 {max(min(M_stray015/sqrt(abs(LsS2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0954 L9TWAXSH03 L2COAXCAB02 {max(min(M_stray015/sqrt(abs(LsS2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0955 L9TWAXSH03 L3COAXCAB02 {max(min(M_stray015/sqrt(abs(LsS2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0956 L9TWAXSH03 L4COAXCAB02 {max(min(M_stray015/sqrt(abs(LsS2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0957 L10TWAXSH03 L1COAXCAB02 {max(min(M_stray015/sqrt(abs(LsS2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0958 L10TWAXSH03 L2COAXCAB02 {max(min(M_stray015/sqrt(abs(LsS2_TWAXSH03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray0959 L10TWAXSH03 L3COAXCAB02 {max(min(M_stray015/sqrt(abs(LsS2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray0960 L10TWAXSH03 L4COAXCAB02 {max(min(M_stray015/sqrt(abs(LsS2_TWAXSH03*LsG2_COAXCAB02)),0.999),-0.999)}
Cstray015 CAPTWAXSH03 n005COAXCAB02 {C_stray015} $ C#005=<C_stray015>
Kstray0961 L1TWAXSH03 L1COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)} $ M#005=<M_stray016>
Kstray0962 L1TWAXSH03 L2COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0963 L1TWAXSH03 L3COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0964 L1TWAXSH03 L4COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0965 L2TWAXSH03 L1COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0966 L2TWAXSH03 L2COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0967 L2TWAXSH03 L3COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0968 L2TWAXSH03 L4COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0969 L3TWAXSH03 L1COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0970 L3TWAXSH03 L2COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0971 L3TWAXSH03 L3COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0972 L3TWAXSH03 L4COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0973 L4TWAXSH03 L1COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0974 L4TWAXSH03 L2COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0975 L4TWAXSH03 L3COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0976 L4TWAXSH03 L4COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0977 L5TWAXSH03 L1COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0978 L5TWAXSH03 L2COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0979 L5TWAXSH03 L3COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0980 L5TWAXSH03 L4COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0981 L6TWAXSH03 L1COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0982 L6TWAXSH03 L2COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0983 L6TWAXSH03 L3COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0984 L6TWAXSH03 L4COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0985 L7TWAXSH03 L1COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0986 L7TWAXSH03 L2COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0987 L7TWAXSH03 L3COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0988 L7TWAXSH03 L4COAXCAB01 {max(min(M_stray016/sqrt(abs(Ls2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0989 L8TWAXSH03 L1COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0990 L8TWAXSH03 L2COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0991 L8TWAXSH03 L3COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0992 L8TWAXSH03 L4COAXCAB01 {max(min(M_stray016/sqrt(abs(LsG2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0993 L9TWAXSH03 L1COAXCAB01 {max(min(M_stray016/sqrt(abs(LsS2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0994 L9TWAXSH03 L2COAXCAB01 {max(min(M_stray016/sqrt(abs(LsS2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0995 L9TWAXSH03 L3COAXCAB01 {max(min(M_stray016/sqrt(abs(LsS2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0996 L9TWAXSH03 L4COAXCAB01 {max(min(M_stray016/sqrt(abs(LsS2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray0997 L10TWAXSH03 L1COAXCAB01 {max(min(M_stray016/sqrt(abs(LsS2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0998 L10TWAXSH03 L2COAXCAB01 {max(min(M_stray016/sqrt(abs(LsS2_TWAXSH03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray0999 L10TWAXSH03 L3COAXCAB01 {max(min(M_stray016/sqrt(abs(LsS2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1000 L10TWAXSH03 L4COAXCAB01 {max(min(M_stray016/sqrt(abs(LsS2_TWAXSH03*LsG2_COAXCAB01)),0.999),-0.999)}
Cstray016 CAPTWAXSH03 n005COAXCAB01 {C_stray016} $ C#005=<C_stray016>
Kstray1001 L1TWAXSH04 L1COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)} $ M#005=<M_stray017>
Kstray1002 L1TWAXSH04 L2COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1003 L1TWAXSH04 L3COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1004 L1TWAXSH04 L4COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1005 L2TWAXSH04 L1COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1006 L2TWAXSH04 L2COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1007 L2TWAXSH04 L3COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1008 L2TWAXSH04 L4COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1009 L3TWAXSH04 L1COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1010 L3TWAXSH04 L2COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1011 L3TWAXSH04 L3COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1012 L3TWAXSH04 L4COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1013 L4TWAXSH04 L1COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1014 L4TWAXSH04 L2COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1015 L4TWAXSH04 L3COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1016 L4TWAXSH04 L4COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1017 L5TWAXSH04 L1COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1018 L5TWAXSH04 L2COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1019 L5TWAXSH04 L3COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1020 L5TWAXSH04 L4COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1021 L6TWAXSH04 L1COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1022 L6TWAXSH04 L2COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1023 L6TWAXSH04 L3COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1024 L6TWAXSH04 L4COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1025 L7TWAXSH04 L1COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1026 L7TWAXSH04 L2COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1027 L7TWAXSH04 L3COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1028 L7TWAXSH04 L4COAXCAB02 {max(min(M_stray017/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1029 L8TWAXSH04 L1COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1030 L8TWAXSH04 L2COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1031 L8TWAXSH04 L3COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1032 L8TWAXSH04 L4COAXCAB02 {max(min(M_stray017/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1033 L9TWAXSH04 L1COAXCAB02 {max(min(M_stray017/sqrt(abs(LsS2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1034 L9TWAXSH04 L2COAXCAB02 {max(min(M_stray017/sqrt(abs(LsS2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1035 L9TWAXSH04 L3COAXCAB02 {max(min(M_stray017/sqrt(abs(LsS2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1036 L9TWAXSH04 L4COAXCAB02 {max(min(M_stray017/sqrt(abs(LsS2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1037 L10TWAXSH04 L1COAXCAB02 {max(min(M_stray017/sqrt(abs(LsS2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1038 L10TWAXSH04 L2COAXCAB02 {max(min(M_stray017/sqrt(abs(LsS2_TWAXSH04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1039 L10TWAXSH04 L3COAXCAB02 {max(min(M_stray017/sqrt(abs(LsS2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1040 L10TWAXSH04 L4COAXCAB02 {max(min(M_stray017/sqrt(abs(LsS2_TWAXSH04*LsG2_COAXCAB02)),0.999),-0.999)}
Cstray017 CAPTWAXSH04 n005COAXCAB02 {C_stray017} $ C#005=<C_stray017>
Kstray1041 L1TWAXSH04 L1COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)} $ M#005=<M_stray018>
Kstray1042 L1TWAXSH04 L2COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1043 L1TWAXSH04 L3COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1044 L1TWAXSH04 L4COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1045 L2TWAXSH04 L1COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1046 L2TWAXSH04 L2COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1047 L2TWAXSH04 L3COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1048 L2TWAXSH04 L4COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1049 L3TWAXSH04 L1COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1050 L3TWAXSH04 L2COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1051 L3TWAXSH04 L3COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1052 L3TWAXSH04 L4COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1053 L4TWAXSH04 L1COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1054 L4TWAXSH04 L2COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1055 L4TWAXSH04 L3COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1056 L4TWAXSH04 L4COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1057 L5TWAXSH04 L1COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1058 L5TWAXSH04 L2COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1059 L5TWAXSH04 L3COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1060 L5TWAXSH04 L4COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1061 L6TWAXSH04 L1COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1062 L6TWAXSH04 L2COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1063 L6TWAXSH04 L3COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1064 L6TWAXSH04 L4COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1065 L7TWAXSH04 L1COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1066 L7TWAXSH04 L2COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1067 L7TWAXSH04 L3COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1068 L7TWAXSH04 L4COAXCAB01 {max(min(M_stray018/sqrt(abs(Ls2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1069 L8TWAXSH04 L1COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1070 L8TWAXSH04 L2COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1071 L8TWAXSH04 L3COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1072 L8TWAXSH04 L4COAXCAB01 {max(min(M_stray018/sqrt(abs(LsG2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1073 L9TWAXSH04 L1COAXCAB01 {max(min(M_stray018/sqrt(abs(LsS2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1074 L9TWAXSH04 L2COAXCAB01 {max(min(M_stray018/sqrt(abs(LsS2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1075 L9TWAXSH04 L3COAXCAB01 {max(min(M_stray018/sqrt(abs(LsS2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1076 L9TWAXSH04 L4COAXCAB01 {max(min(M_stray018/sqrt(abs(LsS2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1077 L10TWAXSH04 L1COAXCAB01 {max(min(M_stray018/sqrt(abs(LsS2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1078 L10TWAXSH04 L2COAXCAB01 {max(min(M_stray018/sqrt(abs(LsS2_TWAXSH04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1079 L10TWAXSH04 L3COAXCAB01 {max(min(M_stray018/sqrt(abs(LsS2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1080 L10TWAXSH04 L4COAXCAB01 {max(min(M_stray018/sqrt(abs(LsS2_TWAXSH04*LsG2_COAXCAB01)),0.999),-0.999)}
Cstray018 CAPTWAXSH04 n005COAXCAB01 {C_stray018} $ C#005=<C_stray018>
Kstray1081 L1COAXCAB03 L1COAXCAB02 {max(min(M_stray019/sqrt(abs(Ls2_COAXCAB03*Ls2_COAXCAB02)),0.999),-0.999)} $ M#005=<M_stray019>
Kstray1082 L1COAXCAB03 L2COAXCAB02 {max(min(M_stray019/sqrt(abs(Ls2_COAXCAB03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1083 L1COAXCAB03 L3COAXCAB02 {max(min(M_stray019/sqrt(abs(Ls2_COAXCAB03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1084 L1COAXCAB03 L4COAXCAB02 {max(min(M_stray019/sqrt(abs(Ls2_COAXCAB03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1085 L2COAXCAB03 L1COAXCAB02 {max(min(M_stray019/sqrt(abs(Ls2_COAXCAB03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1086 L2COAXCAB03 L2COAXCAB02 {max(min(M_stray019/sqrt(abs(Ls2_COAXCAB03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1087 L2COAXCAB03 L3COAXCAB02 {max(min(M_stray019/sqrt(abs(Ls2_COAXCAB03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1088 L2COAXCAB03 L4COAXCAB02 {max(min(M_stray019/sqrt(abs(Ls2_COAXCAB03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1089 L3COAXCAB03 L1COAXCAB02 {max(min(M_stray019/sqrt(abs(LsG2_COAXCAB03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1090 L3COAXCAB03 L2COAXCAB02 {max(min(M_stray019/sqrt(abs(LsG2_COAXCAB03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1091 L3COAXCAB03 L3COAXCAB02 {max(min(M_stray019/sqrt(abs(LsG2_COAXCAB03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1092 L3COAXCAB03 L4COAXCAB02 {max(min(M_stray019/sqrt(abs(LsG2_COAXCAB03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1093 L4COAXCAB03 L1COAXCAB02 {max(min(M_stray019/sqrt(abs(LsG2_COAXCAB03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1094 L4COAXCAB03 L2COAXCAB02 {max(min(M_stray019/sqrt(abs(LsG2_COAXCAB03*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1095 L4COAXCAB03 L3COAXCAB02 {max(min(M_stray019/sqrt(abs(LsG2_COAXCAB03*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1096 L4COAXCAB03 L4COAXCAB02 {max(min(M_stray019/sqrt(abs(LsG2_COAXCAB03*LsG2_COAXCAB02)),0.999),-0.999)}
Cstray019 n005COAXCAB03 n005COAXCAB02 {C_stray019} $ C#005=<C_stray019>
Kstray1097 L1COAXCAB03 L1COAXCAB01 {max(min(M_stray020/sqrt(abs(Ls2_COAXCAB03*Ls2_COAXCAB01)),0.999),-0.999)} $ M#005=<M_stray020>
Kstray1098 L1COAXCAB03 L2COAXCAB01 {max(min(M_stray020/sqrt(abs(Ls2_COAXCAB03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1099 L1COAXCAB03 L3COAXCAB01 {max(min(M_stray020/sqrt(abs(Ls2_COAXCAB03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1100 L1COAXCAB03 L4COAXCAB01 {max(min(M_stray020/sqrt(abs(Ls2_COAXCAB03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1101 L2COAXCAB03 L1COAXCAB01 {max(min(M_stray020/sqrt(abs(Ls2_COAXCAB03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1102 L2COAXCAB03 L2COAXCAB01 {max(min(M_stray020/sqrt(abs(Ls2_COAXCAB03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1103 L2COAXCAB03 L3COAXCAB01 {max(min(M_stray020/sqrt(abs(Ls2_COAXCAB03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1104 L2COAXCAB03 L4COAXCAB01 {max(min(M_stray020/sqrt(abs(Ls2_COAXCAB03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1105 L3COAXCAB03 L1COAXCAB01 {max(min(M_stray020/sqrt(abs(LsG2_COAXCAB03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1106 L3COAXCAB03 L2COAXCAB01 {max(min(M_stray020/sqrt(abs(LsG2_COAXCAB03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1107 L3COAXCAB03 L3COAXCAB01 {max(min(M_stray020/sqrt(abs(LsG2_COAXCAB03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1108 L3COAXCAB03 L4COAXCAB01 {max(min(M_stray020/sqrt(abs(LsG2_COAXCAB03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1109 L4COAXCAB03 L1COAXCAB01 {max(min(M_stray020/sqrt(abs(LsG2_COAXCAB03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1110 L4COAXCAB03 L2COAXCAB01 {max(min(M_stray020/sqrt(abs(LsG2_COAXCAB03*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1111 L4COAXCAB03 L3COAXCAB01 {max(min(M_stray020/sqrt(abs(LsG2_COAXCAB03*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1112 L4COAXCAB03 L4COAXCAB01 {max(min(M_stray020/sqrt(abs(LsG2_COAXCAB03*LsG2_COAXCAB01)),0.999),-0.999)}
Cstray020 n005COAXCAB03 n005COAXCAB01 {C_stray020} $ C#005=<C_stray020>
Kstray1113 L1COAXCAB02 L1COAXCAB01 {max(min(M_stray021/sqrt(abs(Ls2_COAXCAB02*Ls2_COAXCAB01)),0.999),-0.999)} $ M#006=<M_stray021>
Kstray1114 L1COAXCAB02 L2COAXCAB01 {max(min(M_stray021/sqrt(abs(Ls2_COAXCAB02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1115 L1COAXCAB02 L3COAXCAB01 {max(min(M_stray021/sqrt(abs(Ls2_COAXCAB02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1116 L1COAXCAB02 L4COAXCAB01 {max(min(M_stray021/sqrt(abs(Ls2_COAXCAB02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1117 L2COAXCAB02 L1COAXCAB01 {max(min(M_stray021/sqrt(abs(Ls2_COAXCAB02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1118 L2COAXCAB02 L2COAXCAB01 {max(min(M_stray021/sqrt(abs(Ls2_COAXCAB02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1119 L2COAXCAB02 L3COAXCAB01 {max(min(M_stray021/sqrt(abs(Ls2_COAXCAB02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1120 L2COAXCAB02 L4COAXCAB01 {max(min(M_stray021/sqrt(abs(Ls2_COAXCAB02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1121 L3COAXCAB02 L1COAXCAB01 {max(min(M_stray021/sqrt(abs(LsG2_COAXCAB02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1122 L3COAXCAB02 L2COAXCAB01 {max(min(M_stray021/sqrt(abs(LsG2_COAXCAB02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1123 L3COAXCAB02 L3COAXCAB01 {max(min(M_stray021/sqrt(abs(LsG2_COAXCAB02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1124 L3COAXCAB02 L4COAXCAB01 {max(min(M_stray021/sqrt(abs(LsG2_COAXCAB02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1125 L4COAXCAB02 L1COAXCAB01 {max(min(M_stray021/sqrt(abs(LsG2_COAXCAB02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1126 L4COAXCAB02 L2COAXCAB01 {max(min(M_stray021/sqrt(abs(LsG2_COAXCAB02*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1127 L4COAXCAB02 L3COAXCAB01 {max(min(M_stray021/sqrt(abs(LsG2_COAXCAB02*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1128 L4COAXCAB02 L4COAXCAB01 {max(min(M_stray021/sqrt(abs(LsG2_COAXCAB02*LsG2_COAXCAB01)),0.999),-0.999)}
Cstray021 n005COAXCAB02 n005COAXCAB01 {C_stray021} $ C#006=<C_stray021>
Kstray1129 L1COAXCAB04 L1COAXCAB05 {max(min(M_stray022/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB05)),0.999),-0.999)} $ M#007=<M_stray022>
Kstray1130 L1COAXCAB04 L2COAXCAB05 {max(min(M_stray022/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1131 L1COAXCAB04 L3COAXCAB05 {max(min(M_stray022/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1132 L1COAXCAB04 L4COAXCAB05 {max(min(M_stray022/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1133 L2COAXCAB04 L1COAXCAB05 {max(min(M_stray022/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1134 L2COAXCAB04 L2COAXCAB05 {max(min(M_stray022/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1135 L2COAXCAB04 L3COAXCAB05 {max(min(M_stray022/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1136 L2COAXCAB04 L4COAXCAB05 {max(min(M_stray022/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1137 L3COAXCAB04 L1COAXCAB05 {max(min(M_stray022/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1138 L3COAXCAB04 L2COAXCAB05 {max(min(M_stray022/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1139 L3COAXCAB04 L3COAXCAB05 {max(min(M_stray022/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1140 L3COAXCAB04 L4COAXCAB05 {max(min(M_stray022/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1141 L4COAXCAB04 L1COAXCAB05 {max(min(M_stray022/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1142 L4COAXCAB04 L2COAXCAB05 {max(min(M_stray022/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1143 L4COAXCAB04 L3COAXCAB05 {max(min(M_stray022/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1144 L4COAXCAB04 L4COAXCAB05 {max(min(M_stray022/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB05)),0.999),-0.999)}
Cstray022 n005COAXCAB04 n005COAXCAB05 {C_stray022} $ C#007=<C_stray022>
Kstray1145 L1COAXCAB06 L1COAXCAB07 {max(min(M_stray023/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB07)),0.999),-0.999)} $ M#008=<M_stray023>
Kstray1146 L1COAXCAB06 L2COAXCAB07 {max(min(M_stray023/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB07)),0.999),-0.999)}
Kstray1147 L1COAXCAB06 L3COAXCAB07 {max(min(M_stray023/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB07)),0.999),-0.999)}
Kstray1148 L1COAXCAB06 L4COAXCAB07 {max(min(M_stray023/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB07)),0.999),-0.999)}
Kstray1149 L2COAXCAB06 L1COAXCAB07 {max(min(M_stray023/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB07)),0.999),-0.999)}
Kstray1150 L2COAXCAB06 L2COAXCAB07 {max(min(M_stray023/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB07)),0.999),-0.999)}
Kstray1151 L2COAXCAB06 L3COAXCAB07 {max(min(M_stray023/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB07)),0.999),-0.999)}
Kstray1152 L2COAXCAB06 L4COAXCAB07 {max(min(M_stray023/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB07)),0.999),-0.999)}
Kstray1153 L3COAXCAB06 L1COAXCAB07 {max(min(M_stray023/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB07)),0.999),-0.999)}
Kstray1154 L3COAXCAB06 L2COAXCAB07 {max(min(M_stray023/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB07)),0.999),-0.999)}
Kstray1155 L3COAXCAB06 L3COAXCAB07 {max(min(M_stray023/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB07)),0.999),-0.999)}
Kstray1156 L3COAXCAB06 L4COAXCAB07 {max(min(M_stray023/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB07)),0.999),-0.999)}
Kstray1157 L4COAXCAB06 L1COAXCAB07 {max(min(M_stray023/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB07)),0.999),-0.999)}
Kstray1158 L4COAXCAB06 L2COAXCAB07 {max(min(M_stray023/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB07)),0.999),-0.999)}
Kstray1159 L4COAXCAB06 L3COAXCAB07 {max(min(M_stray023/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB07)),0.999),-0.999)}
Kstray1160 L4COAXCAB06 L4COAXCAB07 {max(min(M_stray023/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB07)),0.999),-0.999)}
Cstray023 n005COAXCAB06 n005COAXCAB07 {C_stray023} $ C#008=<C_stray023>
Kstray1161 L1COAXCAB06 L1COAXCAB04 {max(min(M_stray024/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB04)),0.999),-0.999)} $ M#009=<M_stray024>
Kstray1162 L1COAXCAB06 L2COAXCAB04 {max(min(M_stray024/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB04)),0.999),-0.999)}
Kstray1163 L1COAXCAB06 L3COAXCAB04 {max(min(M_stray024/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB04)),0.999),-0.999)}
Kstray1164 L1COAXCAB06 L4COAXCAB04 {max(min(M_stray024/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB04)),0.999),-0.999)}
Kstray1165 L2COAXCAB06 L1COAXCAB04 {max(min(M_stray024/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB04)),0.999),-0.999)}
Kstray1166 L2COAXCAB06 L2COAXCAB04 {max(min(M_stray024/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB04)),0.999),-0.999)}
Kstray1167 L2COAXCAB06 L3COAXCAB04 {max(min(M_stray024/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB04)),0.999),-0.999)}
Kstray1168 L2COAXCAB06 L4COAXCAB04 {max(min(M_stray024/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB04)),0.999),-0.999)}
Kstray1169 L3COAXCAB06 L1COAXCAB04 {max(min(M_stray024/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB04)),0.999),-0.999)}
Kstray1170 L3COAXCAB06 L2COAXCAB04 {max(min(M_stray024/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB04)),0.999),-0.999)}
Kstray1171 L3COAXCAB06 L3COAXCAB04 {max(min(M_stray024/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB04)),0.999),-0.999)}
Kstray1172 L3COAXCAB06 L4COAXCAB04 {max(min(M_stray024/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB04)),0.999),-0.999)}
Kstray1173 L4COAXCAB06 L1COAXCAB04 {max(min(M_stray024/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB04)),0.999),-0.999)}
Kstray1174 L4COAXCAB06 L2COAXCAB04 {max(min(M_stray024/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB04)),0.999),-0.999)}
Kstray1175 L4COAXCAB06 L3COAXCAB04 {max(min(M_stray024/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB04)),0.999),-0.999)}
Kstray1176 L4COAXCAB06 L4COAXCAB04 {max(min(M_stray024/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB04)),0.999),-0.999)}
Cstray024 n005COAXCAB06 n005COAXCAB04 {C_stray024} $ C#009=<C_stray024>
Kstray1177 L1COAXCAB06 L1COAXCAB05 {max(min(M_stray025/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB05)),0.999),-0.999)} $ M#009=<M_stray025>
Kstray1178 L1COAXCAB06 L2COAXCAB05 {max(min(M_stray025/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1179 L1COAXCAB06 L3COAXCAB05 {max(min(M_stray025/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1180 L1COAXCAB06 L4COAXCAB05 {max(min(M_stray025/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1181 L2COAXCAB06 L1COAXCAB05 {max(min(M_stray025/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1182 L2COAXCAB06 L2COAXCAB05 {max(min(M_stray025/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1183 L2COAXCAB06 L3COAXCAB05 {max(min(M_stray025/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1184 L2COAXCAB06 L4COAXCAB05 {max(min(M_stray025/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1185 L3COAXCAB06 L1COAXCAB05 {max(min(M_stray025/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1186 L3COAXCAB06 L2COAXCAB05 {max(min(M_stray025/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1187 L3COAXCAB06 L3COAXCAB05 {max(min(M_stray025/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1188 L3COAXCAB06 L4COAXCAB05 {max(min(M_stray025/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1189 L4COAXCAB06 L1COAXCAB05 {max(min(M_stray025/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1190 L4COAXCAB06 L2COAXCAB05 {max(min(M_stray025/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1191 L4COAXCAB06 L3COAXCAB05 {max(min(M_stray025/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1192 L4COAXCAB06 L4COAXCAB05 {max(min(M_stray025/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB05)),0.999),-0.999)}
Cstray025 n005COAXCAB06 n005COAXCAB05 {C_stray025} $ C#009=<C_stray025>
Kstray1193 L1COAXCAB07 L1COAXCAB04 {max(min(M_stray026/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB04)),0.999),-0.999)} $ M#009=<M_stray026>
Kstray1194 L1COAXCAB07 L2COAXCAB04 {max(min(M_stray026/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB04)),0.999),-0.999)}
Kstray1195 L1COAXCAB07 L3COAXCAB04 {max(min(M_stray026/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB04)),0.999),-0.999)}
Kstray1196 L1COAXCAB07 L4COAXCAB04 {max(min(M_stray026/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB04)),0.999),-0.999)}
Kstray1197 L2COAXCAB07 L1COAXCAB04 {max(min(M_stray026/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB04)),0.999),-0.999)}
Kstray1198 L2COAXCAB07 L2COAXCAB04 {max(min(M_stray026/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB04)),0.999),-0.999)}
Kstray1199 L2COAXCAB07 L3COAXCAB04 {max(min(M_stray026/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB04)),0.999),-0.999)}
Kstray1200 L2COAXCAB07 L4COAXCAB04 {max(min(M_stray026/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB04)),0.999),-0.999)}
Kstray1201 L3COAXCAB07 L1COAXCAB04 {max(min(M_stray026/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB04)),0.999),-0.999)}
Kstray1202 L3COAXCAB07 L2COAXCAB04 {max(min(M_stray026/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB04)),0.999),-0.999)}
Kstray1203 L3COAXCAB07 L3COAXCAB04 {max(min(M_stray026/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB04)),0.999),-0.999)}
Kstray1204 L3COAXCAB07 L4COAXCAB04 {max(min(M_stray026/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB04)),0.999),-0.999)}
Kstray1205 L4COAXCAB07 L1COAXCAB04 {max(min(M_stray026/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB04)),0.999),-0.999)}
Kstray1206 L4COAXCAB07 L2COAXCAB04 {max(min(M_stray026/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB04)),0.999),-0.999)}
Kstray1207 L4COAXCAB07 L3COAXCAB04 {max(min(M_stray026/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB04)),0.999),-0.999)}
Kstray1208 L4COAXCAB07 L4COAXCAB04 {max(min(M_stray026/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB04)),0.999),-0.999)}
Cstray026 n005COAXCAB07 n005COAXCAB04 {C_stray026} $ C#009=<C_stray026>
Kstray1209 L1COAXCAB07 L1COAXCAB05 {max(min(M_stray027/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB05)),0.999),-0.999)} $ M#009=<M_stray027>
Kstray1210 L1COAXCAB07 L2COAXCAB05 {max(min(M_stray027/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1211 L1COAXCAB07 L3COAXCAB05 {max(min(M_stray027/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1212 L1COAXCAB07 L4COAXCAB05 {max(min(M_stray027/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1213 L2COAXCAB07 L1COAXCAB05 {max(min(M_stray027/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1214 L2COAXCAB07 L2COAXCAB05 {max(min(M_stray027/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1215 L2COAXCAB07 L3COAXCAB05 {max(min(M_stray027/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1216 L2COAXCAB07 L4COAXCAB05 {max(min(M_stray027/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1217 L3COAXCAB07 L1COAXCAB05 {max(min(M_stray027/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1218 L3COAXCAB07 L2COAXCAB05 {max(min(M_stray027/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1219 L3COAXCAB07 L3COAXCAB05 {max(min(M_stray027/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1220 L3COAXCAB07 L4COAXCAB05 {max(min(M_stray027/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1221 L4COAXCAB07 L1COAXCAB05 {max(min(M_stray027/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1222 L4COAXCAB07 L2COAXCAB05 {max(min(M_stray027/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB05)),0.999),-0.999)}
Kstray1223 L4COAXCAB07 L3COAXCAB05 {max(min(M_stray027/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB05)),0.999),-0.999)}
Kstray1224 L4COAXCAB07 L4COAXCAB05 {max(min(M_stray027/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB05)),0.999),-0.999)}
Cstray027 n005COAXCAB07 n005COAXCAB05 {C_stray027} $ C#009=<C_stray027>
Kstray1225 L1COAXCAB04 L1TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)} $ M#010=<M_stray028>
Kstray1226 L1COAXCAB04 L2TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1227 L1COAXCAB04 L3TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1228 L1COAXCAB04 L4TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1229 L1COAXCAB04 L5TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1230 L1COAXCAB04 L6TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1231 L1COAXCAB04 L7TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1232 L1COAXCAB04 L8TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1233 L1COAXCAB04 L9TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1234 L1COAXCAB04 L10TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1235 L2COAXCAB04 L1TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1236 L2COAXCAB04 L2TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1237 L2COAXCAB04 L3TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1238 L2COAXCAB04 L4TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1239 L2COAXCAB04 L5TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1240 L2COAXCAB04 L6TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1241 L2COAXCAB04 L7TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1242 L2COAXCAB04 L8TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1243 L2COAXCAB04 L9TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1244 L2COAXCAB04 L10TWAXSH01 {max(min(M_stray028/sqrt(abs(Ls2_COAXCAB04*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1245 L3COAXCAB04 L1TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1246 L3COAXCAB04 L2TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1247 L3COAXCAB04 L3TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1248 L3COAXCAB04 L4TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1249 L3COAXCAB04 L5TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1250 L3COAXCAB04 L6TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1251 L3COAXCAB04 L7TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1252 L3COAXCAB04 L8TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1253 L3COAXCAB04 L9TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1254 L3COAXCAB04 L10TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1255 L4COAXCAB04 L1TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1256 L4COAXCAB04 L2TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1257 L4COAXCAB04 L3TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1258 L4COAXCAB04 L4TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1259 L4COAXCAB04 L5TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1260 L4COAXCAB04 L6TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1261 L4COAXCAB04 L7TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1262 L4COAXCAB04 L8TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1263 L4COAXCAB04 L9TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1264 L4COAXCAB04 L10TWAXSH01 {max(min(M_stray028/sqrt(abs(LsG2_COAXCAB04*LsS2_TWAXSH01)),0.999),-0.999)}
Cstray028 n005COAXCAB04 CAPTWAXSH01 {C_stray028} $ C#010=<C_stray028>
Kstray1265 L1COAXCAB04 L1TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)} $ M#010=<M_stray029>
Kstray1266 L1COAXCAB04 L2TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1267 L1COAXCAB04 L3TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1268 L1COAXCAB04 L4TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1269 L1COAXCAB04 L5TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1270 L1COAXCAB04 L6TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1271 L1COAXCAB04 L7TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1272 L1COAXCAB04 L8TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1273 L1COAXCAB04 L9TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1274 L1COAXCAB04 L10TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1275 L2COAXCAB04 L1TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1276 L2COAXCAB04 L2TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1277 L2COAXCAB04 L3TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1278 L2COAXCAB04 L4TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1279 L2COAXCAB04 L5TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1280 L2COAXCAB04 L6TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1281 L2COAXCAB04 L7TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1282 L2COAXCAB04 L8TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1283 L2COAXCAB04 L9TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1284 L2COAXCAB04 L10TWAXSH02 {max(min(M_stray029/sqrt(abs(Ls2_COAXCAB04*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1285 L3COAXCAB04 L1TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1286 L3COAXCAB04 L2TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1287 L3COAXCAB04 L3TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1288 L3COAXCAB04 L4TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1289 L3COAXCAB04 L5TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1290 L3COAXCAB04 L6TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1291 L3COAXCAB04 L7TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1292 L3COAXCAB04 L8TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1293 L3COAXCAB04 L9TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1294 L3COAXCAB04 L10TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1295 L4COAXCAB04 L1TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1296 L4COAXCAB04 L2TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1297 L4COAXCAB04 L3TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1298 L4COAXCAB04 L4TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1299 L4COAXCAB04 L5TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1300 L4COAXCAB04 L6TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1301 L4COAXCAB04 L7TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1302 L4COAXCAB04 L8TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1303 L4COAXCAB04 L9TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1304 L4COAXCAB04 L10TWAXSH02 {max(min(M_stray029/sqrt(abs(LsG2_COAXCAB04*LsS2_TWAXSH02)),0.999),-0.999)}
Cstray029 n005COAXCAB04 CAPTWAXSH02 {C_stray029} $ C#010=<C_stray029>
Kstray1305 L1COAXCAB04 L1COAXCAB03 {max(min(M_stray030/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB03)),0.999),-0.999)} $ M#010=<M_stray030>
Kstray1306 L1COAXCAB04 L2COAXCAB03 {max(min(M_stray030/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1307 L1COAXCAB04 L3COAXCAB03 {max(min(M_stray030/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1308 L1COAXCAB04 L4COAXCAB03 {max(min(M_stray030/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1309 L2COAXCAB04 L1COAXCAB03 {max(min(M_stray030/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1310 L2COAXCAB04 L2COAXCAB03 {max(min(M_stray030/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1311 L2COAXCAB04 L3COAXCAB03 {max(min(M_stray030/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1312 L2COAXCAB04 L4COAXCAB03 {max(min(M_stray030/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1313 L3COAXCAB04 L1COAXCAB03 {max(min(M_stray030/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1314 L3COAXCAB04 L2COAXCAB03 {max(min(M_stray030/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1315 L3COAXCAB04 L3COAXCAB03 {max(min(M_stray030/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1316 L3COAXCAB04 L4COAXCAB03 {max(min(M_stray030/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1317 L4COAXCAB04 L1COAXCAB03 {max(min(M_stray030/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1318 L4COAXCAB04 L2COAXCAB03 {max(min(M_stray030/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1319 L4COAXCAB04 L3COAXCAB03 {max(min(M_stray030/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1320 L4COAXCAB04 L4COAXCAB03 {max(min(M_stray030/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB03)),0.999),-0.999)}
Cstray030 n005COAXCAB04 n005COAXCAB03 {C_stray030} $ C#010=<C_stray030>
Kstray1321 L1COAXCAB05 L1TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)} $ M#010=<M_stray031>
Kstray1322 L1COAXCAB05 L2TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1323 L1COAXCAB05 L3TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1324 L1COAXCAB05 L4TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1325 L1COAXCAB05 L5TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1326 L1COAXCAB05 L6TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1327 L1COAXCAB05 L7TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1328 L1COAXCAB05 L8TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1329 L1COAXCAB05 L9TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1330 L1COAXCAB05 L10TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1331 L2COAXCAB05 L1TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1332 L2COAXCAB05 L2TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1333 L2COAXCAB05 L3TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1334 L2COAXCAB05 L4TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1335 L2COAXCAB05 L5TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1336 L2COAXCAB05 L6TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1337 L2COAXCAB05 L7TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1338 L2COAXCAB05 L8TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1339 L2COAXCAB05 L9TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1340 L2COAXCAB05 L10TWAXSH01 {max(min(M_stray031/sqrt(abs(Ls2_COAXCAB05*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1341 L3COAXCAB05 L1TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1342 L3COAXCAB05 L2TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1343 L3COAXCAB05 L3TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1344 L3COAXCAB05 L4TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1345 L3COAXCAB05 L5TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1346 L3COAXCAB05 L6TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1347 L3COAXCAB05 L7TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1348 L3COAXCAB05 L8TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1349 L3COAXCAB05 L9TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1350 L3COAXCAB05 L10TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1351 L4COAXCAB05 L1TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1352 L4COAXCAB05 L2TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1353 L4COAXCAB05 L3TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1354 L4COAXCAB05 L4TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1355 L4COAXCAB05 L5TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1356 L4COAXCAB05 L6TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1357 L4COAXCAB05 L7TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1358 L4COAXCAB05 L8TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1359 L4COAXCAB05 L9TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1360 L4COAXCAB05 L10TWAXSH01 {max(min(M_stray031/sqrt(abs(LsG2_COAXCAB05*LsS2_TWAXSH01)),0.999),-0.999)}
Cstray031 n005COAXCAB05 CAPTWAXSH01 {C_stray031} $ C#010=<C_stray031>
Kstray1361 L1COAXCAB05 L1TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)} $ M#010=<M_stray032>
Kstray1362 L1COAXCAB05 L2TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1363 L1COAXCAB05 L3TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1364 L1COAXCAB05 L4TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1365 L1COAXCAB05 L5TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1366 L1COAXCAB05 L6TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1367 L1COAXCAB05 L7TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1368 L1COAXCAB05 L8TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1369 L1COAXCAB05 L9TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1370 L1COAXCAB05 L10TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1371 L2COAXCAB05 L1TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1372 L2COAXCAB05 L2TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1373 L2COAXCAB05 L3TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1374 L2COAXCAB05 L4TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1375 L2COAXCAB05 L5TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1376 L2COAXCAB05 L6TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1377 L2COAXCAB05 L7TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1378 L2COAXCAB05 L8TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1379 L2COAXCAB05 L9TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1380 L2COAXCAB05 L10TWAXSH02 {max(min(M_stray032/sqrt(abs(Ls2_COAXCAB05*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1381 L3COAXCAB05 L1TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1382 L3COAXCAB05 L2TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1383 L3COAXCAB05 L3TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1384 L3COAXCAB05 L4TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1385 L3COAXCAB05 L5TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1386 L3COAXCAB05 L6TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1387 L3COAXCAB05 L7TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1388 L3COAXCAB05 L8TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1389 L3COAXCAB05 L9TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1390 L3COAXCAB05 L10TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1391 L4COAXCAB05 L1TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1392 L4COAXCAB05 L2TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1393 L4COAXCAB05 L3TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1394 L4COAXCAB05 L4TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1395 L4COAXCAB05 L5TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1396 L4COAXCAB05 L6TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1397 L4COAXCAB05 L7TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1398 L4COAXCAB05 L8TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1399 L4COAXCAB05 L9TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1400 L4COAXCAB05 L10TWAXSH02 {max(min(M_stray032/sqrt(abs(LsG2_COAXCAB05*LsS2_TWAXSH02)),0.999),-0.999)}
Cstray032 n005COAXCAB05 CAPTWAXSH02 {C_stray032} $ C#010=<C_stray032>
Kstray1401 L1COAXCAB05 L1COAXCAB03 {max(min(M_stray033/sqrt(abs(Ls2_COAXCAB05*Ls2_COAXCAB03)),0.999),-0.999)} $ M#010=<M_stray033>
Kstray1402 L1COAXCAB05 L2COAXCAB03 {max(min(M_stray033/sqrt(abs(Ls2_COAXCAB05*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1403 L1COAXCAB05 L3COAXCAB03 {max(min(M_stray033/sqrt(abs(Ls2_COAXCAB05*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1404 L1COAXCAB05 L4COAXCAB03 {max(min(M_stray033/sqrt(abs(Ls2_COAXCAB05*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1405 L2COAXCAB05 L1COAXCAB03 {max(min(M_stray033/sqrt(abs(Ls2_COAXCAB05*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1406 L2COAXCAB05 L2COAXCAB03 {max(min(M_stray033/sqrt(abs(Ls2_COAXCAB05*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1407 L2COAXCAB05 L3COAXCAB03 {max(min(M_stray033/sqrt(abs(Ls2_COAXCAB05*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1408 L2COAXCAB05 L4COAXCAB03 {max(min(M_stray033/sqrt(abs(Ls2_COAXCAB05*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1409 L3COAXCAB05 L1COAXCAB03 {max(min(M_stray033/sqrt(abs(LsG2_COAXCAB05*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1410 L3COAXCAB05 L2COAXCAB03 {max(min(M_stray033/sqrt(abs(LsG2_COAXCAB05*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1411 L3COAXCAB05 L3COAXCAB03 {max(min(M_stray033/sqrt(abs(LsG2_COAXCAB05*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1412 L3COAXCAB05 L4COAXCAB03 {max(min(M_stray033/sqrt(abs(LsG2_COAXCAB05*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1413 L4COAXCAB05 L1COAXCAB03 {max(min(M_stray033/sqrt(abs(LsG2_COAXCAB05*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1414 L4COAXCAB05 L2COAXCAB03 {max(min(M_stray033/sqrt(abs(LsG2_COAXCAB05*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1415 L4COAXCAB05 L3COAXCAB03 {max(min(M_stray033/sqrt(abs(LsG2_COAXCAB05*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1416 L4COAXCAB05 L4COAXCAB03 {max(min(M_stray033/sqrt(abs(LsG2_COAXCAB05*LsG2_COAXCAB03)),0.999),-0.999)}
Cstray033 n005COAXCAB05 n005COAXCAB03 {C_stray033} $ C#010=<C_stray033>
Kstray1417 L1COAXCAB06 L1TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)} $ M#011=<M_stray034>
Kstray1418 L1COAXCAB06 L2TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1419 L1COAXCAB06 L3TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1420 L1COAXCAB06 L4TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1421 L1COAXCAB06 L5TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1422 L1COAXCAB06 L6TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1423 L1COAXCAB06 L7TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1424 L1COAXCAB06 L8TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1425 L1COAXCAB06 L9TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1426 L1COAXCAB06 L10TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1427 L2COAXCAB06 L1TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1428 L2COAXCAB06 L2TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1429 L2COAXCAB06 L3TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1430 L2COAXCAB06 L4TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1431 L2COAXCAB06 L5TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1432 L2COAXCAB06 L6TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1433 L2COAXCAB06 L7TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1434 L2COAXCAB06 L8TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1435 L2COAXCAB06 L9TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1436 L2COAXCAB06 L10TWAXSH01 {max(min(M_stray034/sqrt(abs(Ls2_COAXCAB06*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1437 L3COAXCAB06 L1TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1438 L3COAXCAB06 L2TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1439 L3COAXCAB06 L3TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1440 L3COAXCAB06 L4TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1441 L3COAXCAB06 L5TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1442 L3COAXCAB06 L6TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1443 L3COAXCAB06 L7TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1444 L3COAXCAB06 L8TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1445 L3COAXCAB06 L9TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1446 L3COAXCAB06 L10TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1447 L4COAXCAB06 L1TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1448 L4COAXCAB06 L2TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1449 L4COAXCAB06 L3TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1450 L4COAXCAB06 L4TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1451 L4COAXCAB06 L5TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1452 L4COAXCAB06 L6TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1453 L4COAXCAB06 L7TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1454 L4COAXCAB06 L8TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1455 L4COAXCAB06 L9TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1456 L4COAXCAB06 L10TWAXSH01 {max(min(M_stray034/sqrt(abs(LsG2_COAXCAB06*LsS2_TWAXSH01)),0.999),-0.999)}
Cstray034 n005COAXCAB06 CAPTWAXSH01 {C_stray034} $ C#011=<C_stray034>
Kstray1457 L1COAXCAB06 L1TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)} $ M#011=<M_stray035>
Kstray1458 L1COAXCAB06 L2TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1459 L1COAXCAB06 L3TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1460 L1COAXCAB06 L4TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1461 L1COAXCAB06 L5TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1462 L1COAXCAB06 L6TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1463 L1COAXCAB06 L7TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1464 L1COAXCAB06 L8TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1465 L1COAXCAB06 L9TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1466 L1COAXCAB06 L10TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1467 L2COAXCAB06 L1TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1468 L2COAXCAB06 L2TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1469 L2COAXCAB06 L3TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1470 L2COAXCAB06 L4TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1471 L2COAXCAB06 L5TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1472 L2COAXCAB06 L6TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1473 L2COAXCAB06 L7TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1474 L2COAXCAB06 L8TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1475 L2COAXCAB06 L9TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1476 L2COAXCAB06 L10TWAXSH02 {max(min(M_stray035/sqrt(abs(Ls2_COAXCAB06*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1477 L3COAXCAB06 L1TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1478 L3COAXCAB06 L2TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1479 L3COAXCAB06 L3TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1480 L3COAXCAB06 L4TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1481 L3COAXCAB06 L5TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1482 L3COAXCAB06 L6TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1483 L3COAXCAB06 L7TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1484 L3COAXCAB06 L8TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1485 L3COAXCAB06 L9TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1486 L3COAXCAB06 L10TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1487 L4COAXCAB06 L1TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1488 L4COAXCAB06 L2TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1489 L4COAXCAB06 L3TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1490 L4COAXCAB06 L4TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1491 L4COAXCAB06 L5TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1492 L4COAXCAB06 L6TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1493 L4COAXCAB06 L7TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1494 L4COAXCAB06 L8TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1495 L4COAXCAB06 L9TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1496 L4COAXCAB06 L10TWAXSH02 {max(min(M_stray035/sqrt(abs(LsG2_COAXCAB06*LsS2_TWAXSH02)),0.999),-0.999)}
Cstray035 n005COAXCAB06 CAPTWAXSH02 {C_stray035} $ C#011=<C_stray035>
Kstray1497 L1COAXCAB06 L1COAXCAB03 {max(min(M_stray036/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB03)),0.999),-0.999)} $ M#011=<M_stray036>
Kstray1498 L1COAXCAB06 L2COAXCAB03 {max(min(M_stray036/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1499 L1COAXCAB06 L3COAXCAB03 {max(min(M_stray036/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1500 L1COAXCAB06 L4COAXCAB03 {max(min(M_stray036/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1501 L2COAXCAB06 L1COAXCAB03 {max(min(M_stray036/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1502 L2COAXCAB06 L2COAXCAB03 {max(min(M_stray036/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1503 L2COAXCAB06 L3COAXCAB03 {max(min(M_stray036/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1504 L2COAXCAB06 L4COAXCAB03 {max(min(M_stray036/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1505 L3COAXCAB06 L1COAXCAB03 {max(min(M_stray036/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1506 L3COAXCAB06 L2COAXCAB03 {max(min(M_stray036/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1507 L3COAXCAB06 L3COAXCAB03 {max(min(M_stray036/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1508 L3COAXCAB06 L4COAXCAB03 {max(min(M_stray036/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1509 L4COAXCAB06 L1COAXCAB03 {max(min(M_stray036/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1510 L4COAXCAB06 L2COAXCAB03 {max(min(M_stray036/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1511 L4COAXCAB06 L3COAXCAB03 {max(min(M_stray036/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1512 L4COAXCAB06 L4COAXCAB03 {max(min(M_stray036/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB03)),0.999),-0.999)}
Cstray036 n005COAXCAB06 n005COAXCAB03 {C_stray036} $ C#011=<C_stray036>
Kstray1513 L1COAXCAB07 L1TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)} $ M#011=<M_stray037>
Kstray1514 L1COAXCAB07 L2TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1515 L1COAXCAB07 L3TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1516 L1COAXCAB07 L4TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1517 L1COAXCAB07 L5TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1518 L1COAXCAB07 L6TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1519 L1COAXCAB07 L7TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1520 L1COAXCAB07 L8TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1521 L1COAXCAB07 L9TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1522 L1COAXCAB07 L10TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1523 L2COAXCAB07 L1TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1524 L2COAXCAB07 L2TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1525 L2COAXCAB07 L3TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1526 L2COAXCAB07 L4TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1527 L2COAXCAB07 L5TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1528 L2COAXCAB07 L6TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1529 L2COAXCAB07 L7TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1530 L2COAXCAB07 L8TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1531 L2COAXCAB07 L9TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1532 L2COAXCAB07 L10TWAXSH01 {max(min(M_stray037/sqrt(abs(Ls2_COAXCAB07*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1533 L3COAXCAB07 L1TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1534 L3COAXCAB07 L2TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1535 L3COAXCAB07 L3TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1536 L3COAXCAB07 L4TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1537 L3COAXCAB07 L5TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1538 L3COAXCAB07 L6TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1539 L3COAXCAB07 L7TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1540 L3COAXCAB07 L8TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1541 L3COAXCAB07 L9TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1542 L3COAXCAB07 L10TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1543 L4COAXCAB07 L1TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1544 L4COAXCAB07 L2TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1545 L4COAXCAB07 L3TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1546 L4COAXCAB07 L4TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1547 L4COAXCAB07 L5TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1548 L4COAXCAB07 L6TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1549 L4COAXCAB07 L7TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1550 L4COAXCAB07 L8TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1551 L4COAXCAB07 L9TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1552 L4COAXCAB07 L10TWAXSH01 {max(min(M_stray037/sqrt(abs(LsG2_COAXCAB07*LsS2_TWAXSH01)),0.999),-0.999)}
Cstray037 n005COAXCAB07 CAPTWAXSH01 {C_stray037} $ C#011=<C_stray037>
Kstray1553 L1COAXCAB07 L1TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)} $ M#011=<M_stray038>
Kstray1554 L1COAXCAB07 L2TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1555 L1COAXCAB07 L3TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1556 L1COAXCAB07 L4TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1557 L1COAXCAB07 L5TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1558 L1COAXCAB07 L6TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1559 L1COAXCAB07 L7TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1560 L1COAXCAB07 L8TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1561 L1COAXCAB07 L9TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1562 L1COAXCAB07 L10TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1563 L2COAXCAB07 L1TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1564 L2COAXCAB07 L2TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1565 L2COAXCAB07 L3TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1566 L2COAXCAB07 L4TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1567 L2COAXCAB07 L5TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1568 L2COAXCAB07 L6TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1569 L2COAXCAB07 L7TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1570 L2COAXCAB07 L8TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1571 L2COAXCAB07 L9TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1572 L2COAXCAB07 L10TWAXSH02 {max(min(M_stray038/sqrt(abs(Ls2_COAXCAB07*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1573 L3COAXCAB07 L1TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1574 L3COAXCAB07 L2TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1575 L3COAXCAB07 L3TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1576 L3COAXCAB07 L4TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1577 L3COAXCAB07 L5TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1578 L3COAXCAB07 L6TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1579 L3COAXCAB07 L7TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1580 L3COAXCAB07 L8TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1581 L3COAXCAB07 L9TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1582 L3COAXCAB07 L10TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1583 L4COAXCAB07 L1TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1584 L4COAXCAB07 L2TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1585 L4COAXCAB07 L3TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1586 L4COAXCAB07 L4TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1587 L4COAXCAB07 L5TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1588 L4COAXCAB07 L6TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1589 L4COAXCAB07 L7TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1590 L4COAXCAB07 L8TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1591 L4COAXCAB07 L9TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1592 L4COAXCAB07 L10TWAXSH02 {max(min(M_stray038/sqrt(abs(LsG2_COAXCAB07*LsS2_TWAXSH02)),0.999),-0.999)}
Cstray038 n005COAXCAB07 CAPTWAXSH02 {C_stray038} $ C#011=<C_stray038>
Kstray1593 L1COAXCAB07 L1COAXCAB03 {max(min(M_stray039/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB03)),0.999),-0.999)} $ M#011=<M_stray039>
Kstray1594 L1COAXCAB07 L2COAXCAB03 {max(min(M_stray039/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1595 L1COAXCAB07 L3COAXCAB03 {max(min(M_stray039/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1596 L1COAXCAB07 L4COAXCAB03 {max(min(M_stray039/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1597 L2COAXCAB07 L1COAXCAB03 {max(min(M_stray039/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1598 L2COAXCAB07 L2COAXCAB03 {max(min(M_stray039/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1599 L2COAXCAB07 L3COAXCAB03 {max(min(M_stray039/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1600 L2COAXCAB07 L4COAXCAB03 {max(min(M_stray039/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1601 L3COAXCAB07 L1COAXCAB03 {max(min(M_stray039/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1602 L3COAXCAB07 L2COAXCAB03 {max(min(M_stray039/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1603 L3COAXCAB07 L3COAXCAB03 {max(min(M_stray039/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1604 L3COAXCAB07 L4COAXCAB03 {max(min(M_stray039/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1605 L4COAXCAB07 L1COAXCAB03 {max(min(M_stray039/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1606 L4COAXCAB07 L2COAXCAB03 {max(min(M_stray039/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1607 L4COAXCAB07 L3COAXCAB03 {max(min(M_stray039/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1608 L4COAXCAB07 L4COAXCAB03 {max(min(M_stray039/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB03)),0.999),-0.999)}
Cstray039 n005COAXCAB07 n005COAXCAB03 {C_stray039} $ C#011=<C_stray039>
Kstray1609 L1COAXCAB04 L1COAXCAB02 {max(min(M_stray040/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB02)),0.999),-0.999)} $ M#012=<M_stray040>
Kstray1610 L1COAXCAB04 L2COAXCAB02 {max(min(M_stray040/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1611 L1COAXCAB04 L3COAXCAB02 {max(min(M_stray040/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1612 L1COAXCAB04 L4COAXCAB02 {max(min(M_stray040/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1613 L2COAXCAB04 L1COAXCAB02 {max(min(M_stray040/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1614 L2COAXCAB04 L2COAXCAB02 {max(min(M_stray040/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1615 L2COAXCAB04 L3COAXCAB02 {max(min(M_stray040/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1616 L2COAXCAB04 L4COAXCAB02 {max(min(M_stray040/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1617 L3COAXCAB04 L1COAXCAB02 {max(min(M_stray040/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1618 L3COAXCAB04 L2COAXCAB02 {max(min(M_stray040/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1619 L3COAXCAB04 L3COAXCAB02 {max(min(M_stray040/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1620 L3COAXCAB04 L4COAXCAB02 {max(min(M_stray040/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1621 L4COAXCAB04 L1COAXCAB02 {max(min(M_stray040/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1622 L4COAXCAB04 L2COAXCAB02 {max(min(M_stray040/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1623 L4COAXCAB04 L3COAXCAB02 {max(min(M_stray040/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1624 L4COAXCAB04 L4COAXCAB02 {max(min(M_stray040/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB02)),0.999),-0.999)}
Cstray040 n005COAXCAB04 n005COAXCAB02 {C_stray040} $ C#012=<C_stray040>
Kstray1625 L1COAXCAB04 L1COAXCAB01 {max(min(M_stray041/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB01)),0.999),-0.999)} $ M#012=<M_stray041>
Kstray1626 L1COAXCAB04 L2COAXCAB01 {max(min(M_stray041/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1627 L1COAXCAB04 L3COAXCAB01 {max(min(M_stray041/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1628 L1COAXCAB04 L4COAXCAB01 {max(min(M_stray041/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1629 L2COAXCAB04 L1COAXCAB01 {max(min(M_stray041/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1630 L2COAXCAB04 L2COAXCAB01 {max(min(M_stray041/sqrt(abs(Ls2_COAXCAB04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1631 L2COAXCAB04 L3COAXCAB01 {max(min(M_stray041/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1632 L2COAXCAB04 L4COAXCAB01 {max(min(M_stray041/sqrt(abs(Ls2_COAXCAB04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1633 L3COAXCAB04 L1COAXCAB01 {max(min(M_stray041/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1634 L3COAXCAB04 L2COAXCAB01 {max(min(M_stray041/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1635 L3COAXCAB04 L3COAXCAB01 {max(min(M_stray041/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1636 L3COAXCAB04 L4COAXCAB01 {max(min(M_stray041/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1637 L4COAXCAB04 L1COAXCAB01 {max(min(M_stray041/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1638 L4COAXCAB04 L2COAXCAB01 {max(min(M_stray041/sqrt(abs(LsG2_COAXCAB04*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1639 L4COAXCAB04 L3COAXCAB01 {max(min(M_stray041/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1640 L4COAXCAB04 L4COAXCAB01 {max(min(M_stray041/sqrt(abs(LsG2_COAXCAB04*LsG2_COAXCAB01)),0.999),-0.999)}
Cstray041 n005COAXCAB04 n005COAXCAB01 {C_stray041} $ C#012=<C_stray041>
Kstray1641 L1COAXCAB05 L1COAXCAB02 {max(min(M_stray042/sqrt(abs(Ls2_COAXCAB05*Ls2_COAXCAB02)),0.999),-0.999)} $ M#012=<M_stray042>
Kstray1642 L1COAXCAB05 L2COAXCAB02 {max(min(M_stray042/sqrt(abs(Ls2_COAXCAB05*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1643 L1COAXCAB05 L3COAXCAB02 {max(min(M_stray042/sqrt(abs(Ls2_COAXCAB05*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1644 L1COAXCAB05 L4COAXCAB02 {max(min(M_stray042/sqrt(abs(Ls2_COAXCAB05*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1645 L2COAXCAB05 L1COAXCAB02 {max(min(M_stray042/sqrt(abs(Ls2_COAXCAB05*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1646 L2COAXCAB05 L2COAXCAB02 {max(min(M_stray042/sqrt(abs(Ls2_COAXCAB05*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1647 L2COAXCAB05 L3COAXCAB02 {max(min(M_stray042/sqrt(abs(Ls2_COAXCAB05*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1648 L2COAXCAB05 L4COAXCAB02 {max(min(M_stray042/sqrt(abs(Ls2_COAXCAB05*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1649 L3COAXCAB05 L1COAXCAB02 {max(min(M_stray042/sqrt(abs(LsG2_COAXCAB05*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1650 L3COAXCAB05 L2COAXCAB02 {max(min(M_stray042/sqrt(abs(LsG2_COAXCAB05*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1651 L3COAXCAB05 L3COAXCAB02 {max(min(M_stray042/sqrt(abs(LsG2_COAXCAB05*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1652 L3COAXCAB05 L4COAXCAB02 {max(min(M_stray042/sqrt(abs(LsG2_COAXCAB05*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1653 L4COAXCAB05 L1COAXCAB02 {max(min(M_stray042/sqrt(abs(LsG2_COAXCAB05*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1654 L4COAXCAB05 L2COAXCAB02 {max(min(M_stray042/sqrt(abs(LsG2_COAXCAB05*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1655 L4COAXCAB05 L3COAXCAB02 {max(min(M_stray042/sqrt(abs(LsG2_COAXCAB05*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1656 L4COAXCAB05 L4COAXCAB02 {max(min(M_stray042/sqrt(abs(LsG2_COAXCAB05*LsG2_COAXCAB02)),0.999),-0.999)}
Cstray042 n005COAXCAB05 n005COAXCAB02 {C_stray042} $ C#012=<C_stray042>
Kstray1657 L1COAXCAB05 L1COAXCAB01 {max(min(M_stray043/sqrt(abs(Ls2_COAXCAB05*Ls2_COAXCAB01)),0.999),-0.999)} $ M#012=<M_stray043>
Kstray1658 L1COAXCAB05 L2COAXCAB01 {max(min(M_stray043/sqrt(abs(Ls2_COAXCAB05*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1659 L1COAXCAB05 L3COAXCAB01 {max(min(M_stray043/sqrt(abs(Ls2_COAXCAB05*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1660 L1COAXCAB05 L4COAXCAB01 {max(min(M_stray043/sqrt(abs(Ls2_COAXCAB05*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1661 L2COAXCAB05 L1COAXCAB01 {max(min(M_stray043/sqrt(abs(Ls2_COAXCAB05*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1662 L2COAXCAB05 L2COAXCAB01 {max(min(M_stray043/sqrt(abs(Ls2_COAXCAB05*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1663 L2COAXCAB05 L3COAXCAB01 {max(min(M_stray043/sqrt(abs(Ls2_COAXCAB05*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1664 L2COAXCAB05 L4COAXCAB01 {max(min(M_stray043/sqrt(abs(Ls2_COAXCAB05*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1665 L3COAXCAB05 L1COAXCAB01 {max(min(M_stray043/sqrt(abs(LsG2_COAXCAB05*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1666 L3COAXCAB05 L2COAXCAB01 {max(min(M_stray043/sqrt(abs(LsG2_COAXCAB05*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1667 L3COAXCAB05 L3COAXCAB01 {max(min(M_stray043/sqrt(abs(LsG2_COAXCAB05*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1668 L3COAXCAB05 L4COAXCAB01 {max(min(M_stray043/sqrt(abs(LsG2_COAXCAB05*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1669 L4COAXCAB05 L1COAXCAB01 {max(min(M_stray043/sqrt(abs(LsG2_COAXCAB05*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1670 L4COAXCAB05 L2COAXCAB01 {max(min(M_stray043/sqrt(abs(LsG2_COAXCAB05*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1671 L4COAXCAB05 L3COAXCAB01 {max(min(M_stray043/sqrt(abs(LsG2_COAXCAB05*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1672 L4COAXCAB05 L4COAXCAB01 {max(min(M_stray043/sqrt(abs(LsG2_COAXCAB05*LsG2_COAXCAB01)),0.999),-0.999)}
Cstray043 n005COAXCAB05 n005COAXCAB01 {C_stray043} $ C#012=<C_stray043>
Kstray1673 L1COAXCAB06 L1COAXCAB02 {max(min(M_stray044/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB02)),0.999),-0.999)} $ M#013=<M_stray044>
Kstray1674 L1COAXCAB06 L2COAXCAB02 {max(min(M_stray044/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1675 L1COAXCAB06 L3COAXCAB02 {max(min(M_stray044/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1676 L1COAXCAB06 L4COAXCAB02 {max(min(M_stray044/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1677 L2COAXCAB06 L1COAXCAB02 {max(min(M_stray044/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1678 L2COAXCAB06 L2COAXCAB02 {max(min(M_stray044/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1679 L2COAXCAB06 L3COAXCAB02 {max(min(M_stray044/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1680 L2COAXCAB06 L4COAXCAB02 {max(min(M_stray044/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1681 L3COAXCAB06 L1COAXCAB02 {max(min(M_stray044/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1682 L3COAXCAB06 L2COAXCAB02 {max(min(M_stray044/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1683 L3COAXCAB06 L3COAXCAB02 {max(min(M_stray044/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1684 L3COAXCAB06 L4COAXCAB02 {max(min(M_stray044/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1685 L4COAXCAB06 L1COAXCAB02 {max(min(M_stray044/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1686 L4COAXCAB06 L2COAXCAB02 {max(min(M_stray044/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1687 L4COAXCAB06 L3COAXCAB02 {max(min(M_stray044/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1688 L4COAXCAB06 L4COAXCAB02 {max(min(M_stray044/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB02)),0.999),-0.999)}
Cstray044 n005COAXCAB06 n005COAXCAB02 {C_stray044} $ C#013=<C_stray044>
Kstray1689 L1COAXCAB06 L1COAXCAB01 {max(min(M_stray045/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB01)),0.999),-0.999)} $ M#013=<M_stray045>
Kstray1690 L1COAXCAB06 L2COAXCAB01 {max(min(M_stray045/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1691 L1COAXCAB06 L3COAXCAB01 {max(min(M_stray045/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1692 L1COAXCAB06 L4COAXCAB01 {max(min(M_stray045/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1693 L2COAXCAB06 L1COAXCAB01 {max(min(M_stray045/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1694 L2COAXCAB06 L2COAXCAB01 {max(min(M_stray045/sqrt(abs(Ls2_COAXCAB06*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1695 L2COAXCAB06 L3COAXCAB01 {max(min(M_stray045/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1696 L2COAXCAB06 L4COAXCAB01 {max(min(M_stray045/sqrt(abs(Ls2_COAXCAB06*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1697 L3COAXCAB06 L1COAXCAB01 {max(min(M_stray045/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1698 L3COAXCAB06 L2COAXCAB01 {max(min(M_stray045/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1699 L3COAXCAB06 L3COAXCAB01 {max(min(M_stray045/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1700 L3COAXCAB06 L4COAXCAB01 {max(min(M_stray045/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1701 L4COAXCAB06 L1COAXCAB01 {max(min(M_stray045/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1702 L4COAXCAB06 L2COAXCAB01 {max(min(M_stray045/sqrt(abs(LsG2_COAXCAB06*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1703 L4COAXCAB06 L3COAXCAB01 {max(min(M_stray045/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1704 L4COAXCAB06 L4COAXCAB01 {max(min(M_stray045/sqrt(abs(LsG2_COAXCAB06*LsG2_COAXCAB01)),0.999),-0.999)}
Cstray045 n005COAXCAB06 n005COAXCAB01 {C_stray045} $ C#013=<C_stray045>
Kstray1705 L1COAXCAB07 L1COAXCAB02 {max(min(M_stray046/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB02)),0.999),-0.999)} $ M#013=<M_stray046>
Kstray1706 L1COAXCAB07 L2COAXCAB02 {max(min(M_stray046/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1707 L1COAXCAB07 L3COAXCAB02 {max(min(M_stray046/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1708 L1COAXCAB07 L4COAXCAB02 {max(min(M_stray046/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1709 L2COAXCAB07 L1COAXCAB02 {max(min(M_stray046/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1710 L2COAXCAB07 L2COAXCAB02 {max(min(M_stray046/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1711 L2COAXCAB07 L3COAXCAB02 {max(min(M_stray046/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1712 L2COAXCAB07 L4COAXCAB02 {max(min(M_stray046/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1713 L3COAXCAB07 L1COAXCAB02 {max(min(M_stray046/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1714 L3COAXCAB07 L2COAXCAB02 {max(min(M_stray046/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1715 L3COAXCAB07 L3COAXCAB02 {max(min(M_stray046/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1716 L3COAXCAB07 L4COAXCAB02 {max(min(M_stray046/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1717 L4COAXCAB07 L1COAXCAB02 {max(min(M_stray046/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1718 L4COAXCAB07 L2COAXCAB02 {max(min(M_stray046/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1719 L4COAXCAB07 L3COAXCAB02 {max(min(M_stray046/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1720 L4COAXCAB07 L4COAXCAB02 {max(min(M_stray046/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB02)),0.999),-0.999)}
Cstray046 n005COAXCAB07 n005COAXCAB02 {C_stray046} $ C#013=<C_stray046>
Kstray1721 L1COAXCAB07 L1COAXCAB01 {max(min(M_stray047/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB01)),0.999),-0.999)} $ M#013=<M_stray047>
Kstray1722 L1COAXCAB07 L2COAXCAB01 {max(min(M_stray047/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1723 L1COAXCAB07 L3COAXCAB01 {max(min(M_stray047/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1724 L1COAXCAB07 L4COAXCAB01 {max(min(M_stray047/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1725 L2COAXCAB07 L1COAXCAB01 {max(min(M_stray047/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1726 L2COAXCAB07 L2COAXCAB01 {max(min(M_stray047/sqrt(abs(Ls2_COAXCAB07*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1727 L2COAXCAB07 L3COAXCAB01 {max(min(M_stray047/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1728 L2COAXCAB07 L4COAXCAB01 {max(min(M_stray047/sqrt(abs(Ls2_COAXCAB07*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1729 L3COAXCAB07 L1COAXCAB01 {max(min(M_stray047/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1730 L3COAXCAB07 L2COAXCAB01 {max(min(M_stray047/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1731 L3COAXCAB07 L3COAXCAB01 {max(min(M_stray047/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1732 L3COAXCAB07 L4COAXCAB01 {max(min(M_stray047/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1733 L4COAXCAB07 L1COAXCAB01 {max(min(M_stray047/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1734 L4COAXCAB07 L2COAXCAB01 {max(min(M_stray047/sqrt(abs(LsG2_COAXCAB07*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1735 L4COAXCAB07 L3COAXCAB01 {max(min(M_stray047/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1736 L4COAXCAB07 L4COAXCAB01 {max(min(M_stray047/sqrt(abs(LsG2_COAXCAB07*LsG2_COAXCAB01)),0.999),-0.999)}
Cstray047 n005COAXCAB07 n005COAXCAB01 {C_stray047} $ C#013=<C_stray047>
Kstray1737 L1GNDLUG14 L1GNDLUG12 {max(min(M_stray048/sqrt(abs(Rwa1lo*Rwa2lo)),0.999),-0.999)} $ M#014=<M_stray048>
Cstray048 n001GNDLUG14 n001GNDLUG12 {C_stray048} $ C#014=<C_stray048>
Kstray1738 L1GNDLUG14 L1GNDLUG10 {max(min(M_stray049/sqrt(abs(Rwa1lo*Rwa3lo)),0.999),-0.999)} $ M#014=<M_stray049>
Cstray049 n001GNDLUG14 n001GNDLUG10 {C_stray049} $ C#014=<C_stray049>
Kstray1739 L1GNDLUG12 L1GNDLUG10 {max(min(M_stray050/sqrt(abs(Rwa2lo*Rwa3lo)),0.999),-0.999)} $ M#014=<M_stray050>
Cstray050 n001GNDLUG12 n001GNDLUG10 {C_stray050} $ C#014=<C_stray050>
Kstray1740 L1GNDLUG14 L1GNDLUG13 {max(min(M_stray051/sqrt(abs(Rwa1lo*Rwa1hi)),0.999),-0.999)} $ M#015=<M_stray051>
Cstray051 n001GNDLUG14 n001GNDLUG13 {C_stray051} $ C#015=<C_stray051>
Kstray1741 L1GNDLUG14 L1GNDLUG11 {max(min(M_stray052/sqrt(abs(Rwa1lo*Rwa2hi)),0.999),-0.999)} $ M#015=<M_stray052>
Cstray052 n001GNDLUG14 n001GNDLUG11 {C_stray052} $ C#015=<C_stray052>
Kstray1742 L1GNDLUG14 L1GNDLUG09 {max(min(M_stray053/sqrt(abs(Rwa1lo*Rwa3hi)),0.999),-0.999)} $ M#015=<M_stray053>
Cstray053 n001GNDLUG14 n001GNDLUG09 {C_stray053} $ C#015=<C_stray053>
Kstray1743 L1GNDLUG12 L1GNDLUG13 {max(min(M_stray054/sqrt(abs(Rwa2lo*Rwa1hi)),0.999),-0.999)} $ M#015=<M_stray054>
Cstray054 n001GNDLUG12 n001GNDLUG13 {C_stray054} $ C#015=<C_stray054>
Kstray1744 L1GNDLUG12 L1GNDLUG11 {max(min(M_stray055/sqrt(abs(Rwa2lo*Rwa2hi)),0.999),-0.999)} $ M#015=<M_stray055>
Cstray055 n001GNDLUG12 n001GNDLUG11 {C_stray055} $ C#015=<C_stray055>
Kstray1745 L1GNDLUG12 L1GNDLUG09 {max(min(M_stray056/sqrt(abs(Rwa2lo*Rwa3hi)),0.999),-0.999)} $ M#015=<M_stray056>
Cstray056 n001GNDLUG12 n001GNDLUG09 {C_stray056} $ C#015=<C_stray056>
Kstray1746 L1GNDLUG10 L1GNDLUG13 {max(min(M_stray057/sqrt(abs(Rwa3lo*Rwa1hi)),0.999),-0.999)} $ M#015=<M_stray057>
Cstray057 n001GNDLUG10 n001GNDLUG13 {C_stray057} $ C#015=<C_stray057>
Kstray1747 L1GNDLUG10 L1GNDLUG11 {max(min(M_stray058/sqrt(abs(Rwa3lo*Rwa2hi)),0.999),-0.999)} $ M#015=<M_stray058>
Cstray058 n001GNDLUG10 n001GNDLUG11 {C_stray058} $ C#015=<C_stray058>
Kstray1748 L1GNDLUG10 L1GNDLUG09 {max(min(M_stray059/sqrt(abs(Rwa3lo*Rwa3hi)),0.999),-0.999)} $ M#015=<M_stray059>
Cstray059 n001GNDLUG10 n001GNDLUG09 {C_stray059} $ C#015=<C_stray059>
Kstray1749 L1GNDLUG08 L1COAXCAB01 {max(min(M_stray060/sqrt(abs(Lgref*Ls2_COAXCAB01)),0.999),-0.999)} $ M#016=<M_stray060>
Kstray1750 L1GNDLUG08 L2COAXCAB01 {max(min(M_stray060/sqrt(abs(Lgref*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1751 L1GNDLUG08 L3COAXCAB01 {max(min(M_stray060/sqrt(abs(Lgref*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1752 L1GNDLUG08 L4COAXCAB01 {max(min(M_stray060/sqrt(abs(Lgref*LsG2_COAXCAB01)),0.999),-0.999)}
Cstray060 n001GNDLUG08 n005COAXCAB01 {C_stray060} $ C#016=<C_stray060>
Kstray1753 L1GNDLUG08 L1COAXCAB02 {max(min(M_stray061/sqrt(abs(Lgref*Ls2_COAXCAB02)),0.999),-0.999)} $ M#016=<M_stray061>
Kstray1754 L1GNDLUG08 L2COAXCAB02 {max(min(M_stray061/sqrt(abs(Lgref*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1755 L1GNDLUG08 L3COAXCAB02 {max(min(M_stray061/sqrt(abs(Lgref*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1756 L1GNDLUG08 L4COAXCAB02 {max(min(M_stray061/sqrt(abs(Lgref*LsG2_COAXCAB02)),0.999),-0.999)}
Cstray061 n001GNDLUG08 n005COAXCAB02 {C_stray061} $ C#016=<C_stray061>
Kstray1757 L1GNDLUG08 L1COAXCAB03 {max(min(M_stray062/sqrt(abs(Lgref*Ls2_COAXCAB03)),0.999),-0.999)} $ M#016=<M_stray062>
Kstray1758 L1GNDLUG08 L2COAXCAB03 {max(min(M_stray062/sqrt(abs(Lgref*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1759 L1GNDLUG08 L3COAXCAB03 {max(min(M_stray062/sqrt(abs(Lgref*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1760 L1GNDLUG08 L4COAXCAB03 {max(min(M_stray062/sqrt(abs(Lgref*LsG2_COAXCAB03)),0.999),-0.999)}
Cstray062 n001GNDLUG08 n005COAXCAB03 {C_stray062} $ C#016=<C_stray062>
Kstray1761 L1GNDLUG08 L1TWAXSH02 {max(min(M_stray063/sqrt(abs(Lgref*LsG2_TWAXSH02)),0.999),-0.999)} $ M#016=<M_stray063>
Kstray1762 L1GNDLUG08 L2TWAXSH02 {max(min(M_stray063/sqrt(abs(Lgref*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1763 L1GNDLUG08 L3TWAXSH02 {max(min(M_stray063/sqrt(abs(Lgref*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1764 L1GNDLUG08 L4TWAXSH02 {max(min(M_stray063/sqrt(abs(Lgref*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1765 L1GNDLUG08 L5TWAXSH02 {max(min(M_stray063/sqrt(abs(Lgref*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1766 L1GNDLUG08 L6TWAXSH02 {max(min(M_stray063/sqrt(abs(Lgref*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1767 L1GNDLUG08 L7TWAXSH02 {max(min(M_stray063/sqrt(abs(Lgref*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1768 L1GNDLUG08 L8TWAXSH02 {max(min(M_stray063/sqrt(abs(Lgref*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1769 L1GNDLUG08 L9TWAXSH02 {max(min(M_stray063/sqrt(abs(Lgref*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1770 L1GNDLUG08 L10TWAXSH02 {max(min(M_stray063/sqrt(abs(Lgref*LsS2_TWAXSH02)),0.999),-0.999)}
Cstray063 n001GNDLUG08 CAPTWAXSH02 {C_stray063} $ C#016=<C_stray063>
Kstray1771 L1GNDLUG08 L1TWAXSH01 {max(min(M_stray064/sqrt(abs(Lgref*LsG2_TWAXSH01)),0.999),-0.999)} $ M#016=<M_stray064>
Kstray1772 L1GNDLUG08 L2TWAXSH01 {max(min(M_stray064/sqrt(abs(Lgref*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1773 L1GNDLUG08 L3TWAXSH01 {max(min(M_stray064/sqrt(abs(Lgref*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1774 L1GNDLUG08 L4TWAXSH01 {max(min(M_stray064/sqrt(abs(Lgref*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1775 L1GNDLUG08 L5TWAXSH01 {max(min(M_stray064/sqrt(abs(Lgref*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1776 L1GNDLUG08 L6TWAXSH01 {max(min(M_stray064/sqrt(abs(Lgref*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1777 L1GNDLUG08 L7TWAXSH01 {max(min(M_stray064/sqrt(abs(Lgref*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1778 L1GNDLUG08 L8TWAXSH01 {max(min(M_stray064/sqrt(abs(Lgref*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1779 L1GNDLUG08 L9TWAXSH01 {max(min(M_stray064/sqrt(abs(Lgref*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1780 L1GNDLUG08 L10TWAXSH01 {max(min(M_stray064/sqrt(abs(Lgref*LsS2_TWAXSH01)),0.999),-0.999)}
Cstray064 n001GNDLUG08 CAPTWAXSH01 {C_stray064} $ C#016=<C_stray064>
Kstray1781 L1GNDLUG08 L1TWAXSH04 {max(min(M_stray065/sqrt(abs(Lgref*LsG2_TWAXSH04)),0.999),-0.999)} $ M#016=<M_stray065>
Kstray1782 L1GNDLUG08 L2TWAXSH04 {max(min(M_stray065/sqrt(abs(Lgref*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray1783 L1GNDLUG08 L3TWAXSH04 {max(min(M_stray065/sqrt(abs(Lgref*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray1784 L1GNDLUG08 L4TWAXSH04 {max(min(M_stray065/sqrt(abs(Lgref*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray1785 L1GNDLUG08 L5TWAXSH04 {max(min(M_stray065/sqrt(abs(Lgref*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray1786 L1GNDLUG08 L6TWAXSH04 {max(min(M_stray065/sqrt(abs(Lgref*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray1787 L1GNDLUG08 L7TWAXSH04 {max(min(M_stray065/sqrt(abs(Lgref*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray1788 L1GNDLUG08 L8TWAXSH04 {max(min(M_stray065/sqrt(abs(Lgref*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray1789 L1GNDLUG08 L9TWAXSH04 {max(min(M_stray065/sqrt(abs(Lgref*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray1790 L1GNDLUG08 L10TWAXSH04 {max(min(M_stray065/sqrt(abs(Lgref*LsS2_TWAXSH04)),0.999),-0.999)}
Cstray065 n001GNDLUG08 CAPTWAXSH04 {C_stray065} $ C#016=<C_stray065>
Kstray1791 L1GNDLUG08 L1TWAXSH03 {max(min(M_stray066/sqrt(abs(Lgref*LsG2_TWAXSH03)),0.999),-0.999)} $ M#016=<M_stray066>
Kstray1792 L1GNDLUG08 L2TWAXSH03 {max(min(M_stray066/sqrt(abs(Lgref*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray1793 L1GNDLUG08 L3TWAXSH03 {max(min(M_stray066/sqrt(abs(Lgref*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray1794 L1GNDLUG08 L4TWAXSH03 {max(min(M_stray066/sqrt(abs(Lgref*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray1795 L1GNDLUG08 L5TWAXSH03 {max(min(M_stray066/sqrt(abs(Lgref*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray1796 L1GNDLUG08 L6TWAXSH03 {max(min(M_stray066/sqrt(abs(Lgref*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray1797 L1GNDLUG08 L7TWAXSH03 {max(min(M_stray066/sqrt(abs(Lgref*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray1798 L1GNDLUG08 L8TWAXSH03 {max(min(M_stray066/sqrt(abs(Lgref*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray1799 L1GNDLUG08 L9TWAXSH03 {max(min(M_stray066/sqrt(abs(Lgref*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray1800 L1GNDLUG08 L10TWAXSH03 {max(min(M_stray066/sqrt(abs(Lgref*LsS2_TWAXSH03)),0.999),-0.999)}
Cstray066 n001GNDLUG08 CAPTWAXSH03 {C_stray066} $ C#016=<C_stray066>
Kstray1801 L1GNDLUG07 L1COAXCAB01 {max(min(M_stray067/sqrt(abs(Lgrd2*Ls2_COAXCAB01)),0.999),-0.999)} $ M#016=<M_stray067>
Kstray1802 L1GNDLUG07 L2COAXCAB01 {max(min(M_stray067/sqrt(abs(Lgrd2*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1803 L1GNDLUG07 L3COAXCAB01 {max(min(M_stray067/sqrt(abs(Lgrd2*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1804 L1GNDLUG07 L4COAXCAB01 {max(min(M_stray067/sqrt(abs(Lgrd2*LsG2_COAXCAB01)),0.999),-0.999)}
Cstray067 n001GNDLUG07 n005COAXCAB01 {C_stray067} $ C#016=<C_stray067>
Kstray1805 L1GNDLUG07 L1COAXCAB02 {max(min(M_stray068/sqrt(abs(Lgrd2*Ls2_COAXCAB02)),0.999),-0.999)} $ M#016=<M_stray068>
Kstray1806 L1GNDLUG07 L2COAXCAB02 {max(min(M_stray068/sqrt(abs(Lgrd2*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1807 L1GNDLUG07 L3COAXCAB02 {max(min(M_stray068/sqrt(abs(Lgrd2*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1808 L1GNDLUG07 L4COAXCAB02 {max(min(M_stray068/sqrt(abs(Lgrd2*LsG2_COAXCAB02)),0.999),-0.999)}
Cstray068 n001GNDLUG07 n005COAXCAB02 {C_stray068} $ C#016=<C_stray068>
Kstray1809 L1GNDLUG07 L1COAXCAB03 {max(min(M_stray069/sqrt(abs(Lgrd2*Ls2_COAXCAB03)),0.999),-0.999)} $ M#016=<M_stray069>
Kstray1810 L1GNDLUG07 L2COAXCAB03 {max(min(M_stray069/sqrt(abs(Lgrd2*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1811 L1GNDLUG07 L3COAXCAB03 {max(min(M_stray069/sqrt(abs(Lgrd2*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1812 L1GNDLUG07 L4COAXCAB03 {max(min(M_stray069/sqrt(abs(Lgrd2*LsG2_COAXCAB03)),0.999),-0.999)}
Cstray069 n001GNDLUG07 n005COAXCAB03 {C_stray069} $ C#016=<C_stray069>
Kstray1813 L1GNDLUG07 L1TWAXSH02 {max(min(M_stray070/sqrt(abs(Lgrd2*LsG2_TWAXSH02)),0.999),-0.999)} $ M#016=<M_stray070>
Kstray1814 L1GNDLUG07 L2TWAXSH02 {max(min(M_stray070/sqrt(abs(Lgrd2*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1815 L1GNDLUG07 L3TWAXSH02 {max(min(M_stray070/sqrt(abs(Lgrd2*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1816 L1GNDLUG07 L4TWAXSH02 {max(min(M_stray070/sqrt(abs(Lgrd2*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1817 L1GNDLUG07 L5TWAXSH02 {max(min(M_stray070/sqrt(abs(Lgrd2*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1818 L1GNDLUG07 L6TWAXSH02 {max(min(M_stray070/sqrt(abs(Lgrd2*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1819 L1GNDLUG07 L7TWAXSH02 {max(min(M_stray070/sqrt(abs(Lgrd2*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1820 L1GNDLUG07 L8TWAXSH02 {max(min(M_stray070/sqrt(abs(Lgrd2*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1821 L1GNDLUG07 L9TWAXSH02 {max(min(M_stray070/sqrt(abs(Lgrd2*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1822 L1GNDLUG07 L10TWAXSH02 {max(min(M_stray070/sqrt(abs(Lgrd2*LsS2_TWAXSH02)),0.999),-0.999)}
Cstray070 n001GNDLUG07 CAPTWAXSH02 {C_stray070} $ C#016=<C_stray070>
Kstray1823 L1GNDLUG07 L1TWAXSH01 {max(min(M_stray071/sqrt(abs(Lgrd2*LsG2_TWAXSH01)),0.999),-0.999)} $ M#016=<M_stray071>
Kstray1824 L1GNDLUG07 L2TWAXSH01 {max(min(M_stray071/sqrt(abs(Lgrd2*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1825 L1GNDLUG07 L3TWAXSH01 {max(min(M_stray071/sqrt(abs(Lgrd2*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1826 L1GNDLUG07 L4TWAXSH01 {max(min(M_stray071/sqrt(abs(Lgrd2*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1827 L1GNDLUG07 L5TWAXSH01 {max(min(M_stray071/sqrt(abs(Lgrd2*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1828 L1GNDLUG07 L6TWAXSH01 {max(min(M_stray071/sqrt(abs(Lgrd2*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1829 L1GNDLUG07 L7TWAXSH01 {max(min(M_stray071/sqrt(abs(Lgrd2*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1830 L1GNDLUG07 L8TWAXSH01 {max(min(M_stray071/sqrt(abs(Lgrd2*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1831 L1GNDLUG07 L9TWAXSH01 {max(min(M_stray071/sqrt(abs(Lgrd2*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1832 L1GNDLUG07 L10TWAXSH01 {max(min(M_stray071/sqrt(abs(Lgrd2*LsS2_TWAXSH01)),0.999),-0.999)}
Cstray071 n001GNDLUG07 CAPTWAXSH01 {C_stray071} $ C#016=<C_stray071>
Kstray1833 L1GNDLUG07 L1TWAXSH04 {max(min(M_stray072/sqrt(abs(Lgrd2*LsG2_TWAXSH04)),0.999),-0.999)} $ M#016=<M_stray072>
Kstray1834 L1GNDLUG07 L2TWAXSH04 {max(min(M_stray072/sqrt(abs(Lgrd2*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray1835 L1GNDLUG07 L3TWAXSH04 {max(min(M_stray072/sqrt(abs(Lgrd2*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray1836 L1GNDLUG07 L4TWAXSH04 {max(min(M_stray072/sqrt(abs(Lgrd2*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray1837 L1GNDLUG07 L5TWAXSH04 {max(min(M_stray072/sqrt(abs(Lgrd2*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray1838 L1GNDLUG07 L6TWAXSH04 {max(min(M_stray072/sqrt(abs(Lgrd2*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray1839 L1GNDLUG07 L7TWAXSH04 {max(min(M_stray072/sqrt(abs(Lgrd2*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray1840 L1GNDLUG07 L8TWAXSH04 {max(min(M_stray072/sqrt(abs(Lgrd2*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray1841 L1GNDLUG07 L9TWAXSH04 {max(min(M_stray072/sqrt(abs(Lgrd2*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray1842 L1GNDLUG07 L10TWAXSH04 {max(min(M_stray072/sqrt(abs(Lgrd2*LsS2_TWAXSH04)),0.999),-0.999)}
Cstray072 n001GNDLUG07 CAPTWAXSH04 {C_stray072} $ C#016=<C_stray072>
Kstray1843 L1GNDLUG07 L1TWAXSH03 {max(min(M_stray073/sqrt(abs(Lgrd2*LsG2_TWAXSH03)),0.999),-0.999)} $ M#016=<M_stray073>
Kstray1844 L1GNDLUG07 L2TWAXSH03 {max(min(M_stray073/sqrt(abs(Lgrd2*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray1845 L1GNDLUG07 L3TWAXSH03 {max(min(M_stray073/sqrt(abs(Lgrd2*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray1846 L1GNDLUG07 L4TWAXSH03 {max(min(M_stray073/sqrt(abs(Lgrd2*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray1847 L1GNDLUG07 L5TWAXSH03 {max(min(M_stray073/sqrt(abs(Lgrd2*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray1848 L1GNDLUG07 L6TWAXSH03 {max(min(M_stray073/sqrt(abs(Lgrd2*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray1849 L1GNDLUG07 L7TWAXSH03 {max(min(M_stray073/sqrt(abs(Lgrd2*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray1850 L1GNDLUG07 L8TWAXSH03 {max(min(M_stray073/sqrt(abs(Lgrd2*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray1851 L1GNDLUG07 L9TWAXSH03 {max(min(M_stray073/sqrt(abs(Lgrd2*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray1852 L1GNDLUG07 L10TWAXSH03 {max(min(M_stray073/sqrt(abs(Lgrd2*LsS2_TWAXSH03)),0.999),-0.999)}
Cstray073 n001GNDLUG07 CAPTWAXSH03 {C_stray073} $ C#016=<C_stray073>
Kstray1853 L1GNDLUG03 L1COAXCAB01 {max(min(M_stray074/sqrt(abs(Lsrc*Ls2_COAXCAB01)),0.999),-0.999)} $ M#016=<M_stray074>
Kstray1854 L1GNDLUG03 L2COAXCAB01 {max(min(M_stray074/sqrt(abs(Lsrc*Ls2_COAXCAB01)),0.999),-0.999)}
Kstray1855 L1GNDLUG03 L3COAXCAB01 {max(min(M_stray074/sqrt(abs(Lsrc*LsG2_COAXCAB01)),0.999),-0.999)}
Kstray1856 L1GNDLUG03 L4COAXCAB01 {max(min(M_stray074/sqrt(abs(Lsrc*LsG2_COAXCAB01)),0.999),-0.999)}
Cstray074 n001GNDLUG03 n005COAXCAB01 {C_stray074} $ C#016=<C_stray074>
Kstray1857 L1GNDLUG03 L1COAXCAB02 {max(min(M_stray075/sqrt(abs(Lsrc*Ls2_COAXCAB02)),0.999),-0.999)} $ M#016=<M_stray075>
Kstray1858 L1GNDLUG03 L2COAXCAB02 {max(min(M_stray075/sqrt(abs(Lsrc*Ls2_COAXCAB02)),0.999),-0.999)}
Kstray1859 L1GNDLUG03 L3COAXCAB02 {max(min(M_stray075/sqrt(abs(Lsrc*LsG2_COAXCAB02)),0.999),-0.999)}
Kstray1860 L1GNDLUG03 L4COAXCAB02 {max(min(M_stray075/sqrt(abs(Lsrc*LsG2_COAXCAB02)),0.999),-0.999)}
Cstray075 n001GNDLUG03 n005COAXCAB02 {C_stray075} $ C#016=<C_stray075>
Kstray1861 L1GNDLUG03 L1COAXCAB03 {max(min(M_stray076/sqrt(abs(Lsrc*Ls2_COAXCAB03)),0.999),-0.999)} $ M#016=<M_stray076>
Kstray1862 L1GNDLUG03 L2COAXCAB03 {max(min(M_stray076/sqrt(abs(Lsrc*Ls2_COAXCAB03)),0.999),-0.999)}
Kstray1863 L1GNDLUG03 L3COAXCAB03 {max(min(M_stray076/sqrt(abs(Lsrc*LsG2_COAXCAB03)),0.999),-0.999)}
Kstray1864 L1GNDLUG03 L4COAXCAB03 {max(min(M_stray076/sqrt(abs(Lsrc*LsG2_COAXCAB03)),0.999),-0.999)}
Cstray076 n001GNDLUG03 n005COAXCAB03 {C_stray076} $ C#016=<C_stray076>
Kstray1865 L1GNDLUG03 L1TWAXSH02 {max(min(M_stray077/sqrt(abs(Lsrc*LsG2_TWAXSH02)),0.999),-0.999)} $ M#016=<M_stray077>
Kstray1866 L1GNDLUG03 L2TWAXSH02 {max(min(M_stray077/sqrt(abs(Lsrc*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1867 L1GNDLUG03 L3TWAXSH02 {max(min(M_stray077/sqrt(abs(Lsrc*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1868 L1GNDLUG03 L4TWAXSH02 {max(min(M_stray077/sqrt(abs(Lsrc*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1869 L1GNDLUG03 L5TWAXSH02 {max(min(M_stray077/sqrt(abs(Lsrc*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1870 L1GNDLUG03 L6TWAXSH02 {max(min(M_stray077/sqrt(abs(Lsrc*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1871 L1GNDLUG03 L7TWAXSH02 {max(min(M_stray077/sqrt(abs(Lsrc*Ls2_TWAXSH02)),0.999),-0.999)}
Kstray1872 L1GNDLUG03 L8TWAXSH02 {max(min(M_stray077/sqrt(abs(Lsrc*LsG2_TWAXSH02)),0.999),-0.999)}
Kstray1873 L1GNDLUG03 L9TWAXSH02 {max(min(M_stray077/sqrt(abs(Lsrc*LsS2_TWAXSH02)),0.999),-0.999)}
Kstray1874 L1GNDLUG03 L10TWAXSH02 {max(min(M_stray077/sqrt(abs(Lsrc*LsS2_TWAXSH02)),0.999),-0.999)}
Cstray077 n001GNDLUG03 CAPTWAXSH02 {C_stray077} $ C#016=<C_stray077>
Kstray1875 L1GNDLUG03 L1TWAXSH01 {max(min(M_stray078/sqrt(abs(Lsrc*LsG2_TWAXSH01)),0.999),-0.999)} $ M#016=<M_stray078>
Kstray1876 L1GNDLUG03 L2TWAXSH01 {max(min(M_stray078/sqrt(abs(Lsrc*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1877 L1GNDLUG03 L3TWAXSH01 {max(min(M_stray078/sqrt(abs(Lsrc*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1878 L1GNDLUG03 L4TWAXSH01 {max(min(M_stray078/sqrt(abs(Lsrc*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1879 L1GNDLUG03 L5TWAXSH01 {max(min(M_stray078/sqrt(abs(Lsrc*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1880 L1GNDLUG03 L6TWAXSH01 {max(min(M_stray078/sqrt(abs(Lsrc*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1881 L1GNDLUG03 L7TWAXSH01 {max(min(M_stray078/sqrt(abs(Lsrc*Ls2_TWAXSH01)),0.999),-0.999)}
Kstray1882 L1GNDLUG03 L8TWAXSH01 {max(min(M_stray078/sqrt(abs(Lsrc*LsG2_TWAXSH01)),0.999),-0.999)}
Kstray1883 L1GNDLUG03 L9TWAXSH01 {max(min(M_stray078/sqrt(abs(Lsrc*LsS2_TWAXSH01)),0.999),-0.999)}
Kstray1884 L1GNDLUG03 L10TWAXSH01 {max(min(M_stray078/sqrt(abs(Lsrc*LsS2_TWAXSH01)),0.999),-0.999)}
Cstray078 n001GNDLUG03 CAPTWAXSH01 {C_stray078} $ C#016=<C_stray078>
Kstray1885 L1GNDLUG03 L1TWAXSH04 {max(min(M_stray079/sqrt(abs(Lsrc*LsG2_TWAXSH04)),0.999),-0.999)} $ M#016=<M_stray079>
Kstray1886 L1GNDLUG03 L2TWAXSH04 {max(min(M_stray079/sqrt(abs(Lsrc*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray1887 L1GNDLUG03 L3TWAXSH04 {max(min(M_stray079/sqrt(abs(Lsrc*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray1888 L1GNDLUG03 L4TWAXSH04 {max(min(M_stray079/sqrt(abs(Lsrc*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray1889 L1GNDLUG03 L5TWAXSH04 {max(min(M_stray079/sqrt(abs(Lsrc*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray1890 L1GNDLUG03 L6TWAXSH04 {max(min(M_stray079/sqrt(abs(Lsrc*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray1891 L1GNDLUG03 L7TWAXSH04 {max(min(M_stray079/sqrt(abs(Lsrc*Ls2_TWAXSH04)),0.999),-0.999)}
Kstray1892 L1GNDLUG03 L8TWAXSH04 {max(min(M_stray079/sqrt(abs(Lsrc*LsG2_TWAXSH04)),0.999),-0.999)}
Kstray1893 L1GNDLUG03 L9TWAXSH04 {max(min(M_stray079/sqrt(abs(Lsrc*LsS2_TWAXSH04)),0.999),-0.999)}
Kstray1894 L1GNDLUG03 L10TWAXSH04 {max(min(M_stray079/sqrt(abs(Lsrc*LsS2_TWAXSH04)),0.999),-0.999)}
Cstray079 n001GNDLUG03 CAPTWAXSH04 {C_stray079} $ C#016=<C_stray079>
Kstray1895 L1GNDLUG03 L1TWAXSH03 {max(min(M_stray080/sqrt(abs(Lsrc*LsG2_TWAXSH03)),0.999),-0.999)} $ M#016=<M_stray080>
Kstray1896 L1GNDLUG03 L2TWAXSH03 {max(min(M_stray080/sqrt(abs(Lsrc*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray1897 L1GNDLUG03 L3TWAXSH03 {max(min(M_stray080/sqrt(abs(Lsrc*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray1898 L1GNDLUG03 L4TWAXSH03 {max(min(M_stray080/sqrt(abs(Lsrc*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray1899 L1GNDLUG03 L5TWAXSH03 {max(min(M_stray080/sqrt(abs(Lsrc*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray1900 L1GNDLUG03 L6TWAXSH03 {max(min(M_stray080/sqrt(abs(Lsrc*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray1901 L1GNDLUG03 L7TWAXSH03 {max(min(M_stray080/sqrt(abs(Lsrc*Ls2_TWAXSH03)),0.999),-0.999)}
Kstray1902 L1GNDLUG03 L8TWAXSH03 {max(min(M_stray080/sqrt(abs(Lsrc*LsG2_TWAXSH03)),0.999),-0.999)}
Kstray1903 L1GNDLUG03 L9TWAXSH03 {max(min(M_stray080/sqrt(abs(Lsrc*LsS2_TWAXSH03)),0.999),-0.999)}
Kstray1904 L1GNDLUG03 L10TWAXSH03 {max(min(M_stray080/sqrt(abs(Lsrc*LsS2_TWAXSH03)),0.999),-0.999)}
Cstray080 n001GNDLUG03 CAPTWAXSH03 {C_stray080} $ C#016=<C_stray080>

.end

